`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OA2cDxxBBgQGJMp2pxvIcb9dg8Uqwmv+0eyEdSECDu3UgdHiXU5FeBOB2Q9h9uII0FkFHF8ZM/p5
QCk1gyZuNA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ohw3/ONQPF4YSQ9T4UlhV3QIxoCPQR4nSH8nk5PkpXa2YESP9l5Ukzz3ov2c4s0uNC7340gxwGIh
iZiO71DkVAEONuxBbBoBIz9wl8KBcu3gIWYM3qoATzEBCvJUsWW3y7x4irWQVePt8OSzl7ugyAKH
Gavs/n2UAAo3JGr9nuQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qbQdmKpXGCQroM/9Mx26/oA5UfkaVHlnKnkEDXAiffyr+pAS4Xq2B/0/lqmbCYBBKnZpRSPoWUEs
Cg1/IqWvWntatpU9JwJ+hjvSRkztujxk9id6jXnKk8AFHe+y36LqoKhVdARle9zcy0G4UlY4ScPP
z18tJGZn1cVPNUr3wbHIKRZS/pdZdBjPIkpZzfpmtwAPWyBT4InH2oT1IUVra4E4Lbc2JeIXcpQI
MA4GDr2IGv/Enl3BKXEt0JzX1tZtq1bzklY6XMcUl1o97QwbFOZa1aUWgVBRRA1AJNIiMyg5Pvfc
Q9phtLshsSkW42KhxQMiXf2l/0OZGMvjsliZOA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ch1JwuARongvYA6wwxtZ9HrijShX8v/T8gJft+KazH/83xQ8WQuf2Auf0DEkLYqXb6lmqjTo5Qv3
/UW4me8gr16uhQcbbM5vhT7Yrb0J0W1xruMlQiO2JNDG9r1RQx2OSK1yi0pPBLLOAlVkKSsgWZbS
tIQhtAj4DXc1oOc5vjpuzgyZ5MsedeXKnOkmG8dO+YW3o63NkPAu9Pl4lAB7oGQEnvua9zRMAsi0
edkVgJdX2DsBhIkBrWZRXQ3TUKGFyrcemkBYBAN/p3IwcmqxU8VD8smJrfUw5ftrr5164WnARz6x
2zZZlLCtzlHvT3Onbva+EKM3a4AioOcXu6Kjag==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VT7lyAYu7/weMOfLvOM+SHZmAAVV6GMaD3gr7ZSNU8JfV9HIoUTxp6J0mJdeOKs3tYYlqi6cF+Qo
F8YCUKXluoy1gcptygDK7q//Xh7zBwLcSKdoUJr/Arnk4ijKQuEZ9JjH98tsD1GIA6B0EUQRclHC
FwSksULSbpayYa7tjvYuijf3sJDtJFxV+GTeKDKTRe8W0jHosQUN+0aKY8WRP/nt7ccDxmn0IZyv
NYwNf0lrWjEC4Ki1WiMukH+NDrbYZZ4V7XSuq11etS2vz0dQpM0oVQxT3DWkod7qrSaHvHyK9moY
KzDcXWkyU3VpqGrxPWl9DJP6lEv2rVhdkpjMbA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XgmFRGaDq2b3xpHvzH+IwGP/IQNDsWlcao685okhs0AfoeD4RtvYCy+nfvG7Y5DWm1xA4Wa046Ju
gEBXPOzaNoAltTfF+odHBTEi+5zMk9gbAJjMmAmBq1RIDStwIFRdEfdyaG+BfFkpmz+MiAGgdUn2
avVOBrCw9WUXA0b+vy0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pjB2Cz+0cSVKp4du1DXMN5l66IUTXx3HaY0OfcBMe+msmACV9SKLQqpbiwy2Glq6Nzrvx960qHGd
FjDXHMKbGPzR33ri6HWVEvLoTZbPfVkX6Jn/yPiNAUbCYBZ6kq0pXUAH3rpN1nE+Eg0wUdWaE9dJ
46214wdWThgp/a2oUEhsBDNuz850Vvo9f3HJGHeUizN/IviKOQCBxQstk1qRDYXVGyiW/vtBTPCL
wVJAZ1C0anyhQAS40N1AKpX8bV9joriwf9jvkmWmBSZB/t12s9UVHmf4Wjyk3vJ2u5s5QKMwb1ag
7LyWm/+cXV1dKHMIaYTLYX6X86whqonJjzSw6g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 261312)
`protect data_block
NcJciS9TpdEiLy7CQ42EdoB4M5rErP0yymQ7zO9/G7AlX9x+FBB5gQxwcNZuRnlBagFWN1+y/kPp
tZx4LLbVA7MReIaHCN1isTK4ijYaAxrJguG8w9B0/vjQmfJl4F4iIbF2c/CWxn4VYr4M0kWhL/Ts
JykLF2g+qKNCxJGQv3yKwXrdgp7a+MzDfpaAR1Pk46i0V3AZZGUZmK9nqWc0w5PHauDHc1O+EK9V
zNzyiRc/A0QEWQ3/izn++cFHjmxMBbYKeNx6iWvuPdYTk42qpeKeIA84xZ1ADk8+H0SQftXBFvnt
HpIpTO54GyKoA3uZb/d7d19jKzG5V7kcp9LkhTeq+CMPKjskhohPxIyILDt4UA7AzSpGG3xdn8ND
g+Qi9l7F+GMtITKhKNa2yuBL4kIG+lOiqd9rVSEZzREkjMbnzWAoqPJRUZ+qfILCbHQPINDHQ946
GuN+Vc9y0w6YK9iwOW3FltEuQyvopk/IIGGqIVLMzHjEfmlxkVLqjVOrUdzYSPeHtXY7Ex0gTNe9
3iVosTFh0NDZz0ilrJ+rfqKHQ+QtlgZtm0LIIAE0IeQsRACEnjSMLysXXuRDMBxe6/tmqvzFaknr
ILlfmzXg8987VwUFaBvzbmTFOQ+A9MtsjtAERv0hI+W/W+IHyiyJPJv3RCoJGnNleWSkH8aXxoQ/
+c+Tao5wH0RszzipxwTfgOhrcgC8pQNxHOmDfNaNC7Knire/hZD+YZx8vuaw+/6EDCSLUSTOEhZB
eyPGqNU9cG9XbSLT4slv1NlFOEYbEKRMr5r9tbtkKfx4DbClQDnksS7bZvNtQspy24BuOdFqhGlb
b8sWW07VsOoMaC1qgsxY3h5yuoQqf1Lmxdu5tES+D6dvYlWYTV4kG7Hhiqj62qovgrUFgEi74JuH
kFmZLREaG90uDpVubNUjmxC7lsTRV0m/aHli8uSVLyXvndvmdF7AHBcU7n+k3WjK/1hNxAZqjmkE
Ch6S0kKsGcbNwxgf3WSbkXqSRA9q2wBGrgk32IKKYJa531pij6IDcT9R8WDvf/MWq5EX5GYRVBZe
Yfb+gPdxmXRRxgLlte37zAk6s02p8BNxZOZKXBbmvp5jwlT2nZfnWtIbyJQMsBhZh4/2RHYXYev/
MnzrjhVum3IrrGpFt8Ihma41C5eIiqMYClDyaTP38zXyMrx1XgTgwdKccafwiejL6It3TEsSOZzP
EhyMXkWdrQPAkX2zCalLcbsSsw3nSDtinzelciLRq3wViD4YhioJ5H4ZP4iQyoT4NhGoQFaV0BB2
KZLbILm4kb0FqjVWCGPiJlUYjERHfu3NqX1JxP/fYfta3Uvqb76NQfoNWGtkQ9PDGgNGkre9DNvp
Hnxm09FxTNHl2Y4mRvB8Te15UulnbbLR+WKUUT9SBVE6oJ08qMqcmkBAwsPRrepz564KzaVd/Ugu
Zwx5OwJD/G+8G7ckL8pnhkBxucz+A1+0R3ntT+ZGGuPSh/XnAZ2i33bOUX5ZwqV0ZZYdOJojd4NR
q5+5SExT1SN/wXnTT0FEJc2ysTbLjDVS3KIwonzTUUycUhmvpvzOkmkcAIW8fE+Kj9H7b3vxH3kw
uy2Nj6wobuqMjCDviXM0rpanOqIgKgfnkPxfXMaFzCny31xL1Ey2haVmM2Ual1zROXL6qtx85qBC
C0fgTA6VDdRyKYmD2k3jElXOkMJ6LkNPI5OHdbRNVgYRibTAI8Qhuq6z1h76EXRaYtxDlHZ191P6
FnUrVeUqIhwk6rb6eBk/iv/56nOx7OE/vExI8kRgPG/ZSeyebpY/VrgVJBVfKmI2Ug0YH6XBRM2C
okDOpTvAJo3XQwdC0rtf83pavnUcHcUPVPQQ8gsQPtJCXQYQ7nhUMRtO6zMTp9Be1y48fi4RUssk
8luWdND6UQ4tcpOv4gzoRafimgtehHofvZNu6CmJzWWPRVAu8dOBpKFKif4i7yVYNyKKlO0Lat1l
Z997/OHHhXiNf/+MCrCr5N35nPzQm/HYVS2drRgaiShygmxQNp6TCFMN1vOTT8sDvLX4obimM8+b
TJ8WDeTMf4hoz9bhd/693O1rI27sdrvtbDKCBRUCouG7/lts7abz3YGRsfGgm5HRsUJVGl0nt+Gg
3tVrUrO9R2PG4QUUSWr14eD4GM3qNqnrqmrXTMmFf/Q7oOocqE9dwKfVYm/Nm7HvLxclbeAmGxDU
26ohtdB+ivoUYraALmnecBvUChU7fVGH6/wotQ9nwgWq8rFsrWJSqiDuA3IO1aE64SuiWXLT2rs7
vXak+UoaHacxzcR+JcS3DlMrC+fILkNQTHu2/8EdqtobNduL0y05r6cePTJefJWn3sYzO2273MLk
c7hutrzQ0ruv/wKktZbTxkl9yQ8/b0tsiFWXYzSL9rqPtUijZd/64sRWxmnX7ESsj5Fa0rQ1rYZi
/cG8PvCp3agTR3XR00jvvz6mPXCn784WJO4axiS+9iWe1DDVNGfcCrWn2WwWOB+wVqPzZrWDrUQy
hiWkTkms7Qm3iN/V50cYfkzjIx9NHZXaLQo8vU26JRnv4+hEaE9xSBbGGilgqO+ikfpA+CPEEZSj
WIucf5XNUGi3Sf5RENQQ2Rklz79/6v87DT+t2uc3YKZujXtwBUOkDEpiDRT5Ghl5T4ReP4zEW4fC
NQ9yTvW0vgF2OfF4XZ6GLZ/0td6PoCCSKvCNccA1dPeAX9Qy5TirFfzFAxooDyWU31XiiyU7sau4
xsIYiRf/eGr+2U/eAj6DP7HHBnsY2s1zf28koDuVkd5WAmWFb2YQqdw/XGfuetEafpJPtRg4q7HO
rZb68/AtFdFIQ2jY0HpguUpYhoGJueNXeqhs/LdLlarpdeQJqaMKrKOaYRvgN+mjoLGw6yLyzOvt
FWeUyXvfPR6+9ixqnspuNktxHrxr3tG05c6oH3/m+CWMtHQjy1tTZNunYBleM2c+nKIxhoV/V4FW
WyNTTdV0j290ET6nRguYqV16uy0II8Mc/Ov0oapgoYKqZIqsSA8rOoC2lKyPUhj+k9/J593YGqhr
dPa4ldB6Fm2jpgu0rTs9gawm0AZyLLo+RKRazJH+QmbwFBb3Cs+s8CEsvG0ylSac3DPze1dNHRy2
BBYxuXOgzLW3jsYmqioqgYBOoKmvvTni/j0foeg0tWM7koLzAREEiMer7eID1liYhlR9rO4bpQTT
BN937ZSj4e4JyVtL2zmHE7c+Kc6Vl5MSIwC7doSlNFYHUs+j37Eqx1fBswAiKlkoDD83W8DzG6ED
raV2HAJNuUKAT/nT1wQDmNzlD4qejk9S+6PuK8ARsOc0vltbx1a9bB1/CXtzsQjVj6cIUpoHQx2z
09EaE/u9jfBUmUY9mC6sQfGgSddBZyX2flImJ5Xrc36odhChsIiKlMxdhXUrVunDnYO5vuCZh98o
mLQWRkDpOu6TicQBQYQZZf04c0UqtLl0ww/3q7jpSwsHrIokFTw531xuoLs8XbmMjy5hEpSAW4dp
qS636AKcAafb9mWUynA43bhWaO8ZOpPkIYZvTO7ncvFkSc/TmljCeznMIrW7emEYuYENBCZUTckW
lqEcdnKInrzU085i2uf+0FBKTeI5REa6NgDN1PK7q5Hcjm31Wv/iTHhKA5mIpye95uhOZZq+8EzQ
xM92/HS8hbA++lNTAppHDaXw/a0ArTmVTRaFs25VYQ0ZvWNYlxwWVbktIvCM36f95QVMQ4SLAQgK
FgZXPJTWeY9XU+J4BIwrocBKRXUb8+3TLqncZQzqcueE8XAg2aJz7YVfubRYGPRsZLT9gOMuAPeB
7THOUYCYqXuHNs2oo+ozpAnjY4FhyympYQGuPkWVzDUyDQlM2P+rgqTMvBwXEntXHEHJaItDTke5
qgrDJHq7obv2msgx1T9GZhn0EkjUm3WaVJeJ4A6VPYPk/42FlqGRh6XYjDuxnizGNxWm2Uz5JXM2
Vamy/qbRS0LUzfj12x7heDqM7/WjaaIlUvyojiGI8QQahBaMzj1UdTW4gdOU6lrVW0pUIwzQkx1o
vf9iSLJbOt+sV9XtT7bc28h13f59mMGB4Y+oafNE103oWeWZZ3GhPutYaVpuwiex/5fiIa4phqaQ
+8MTitDf8YEjm97iio2dHIR0fG8uLb50/65Kvhlinvc1n7xajHFu7lL6mi5ZXLq6MqkULv1ioPxq
TIwUFzvjkgsbBY9VtLH1ue+1n/k8qCO3lNKXdYdhjk7HH87o64ZVTKOrjoYbwnCaFyFgqTTNc3T/
1uQMzIJGlc/X9sbK5AXnzoKgTB9USFrqYeF0nN1m2Tcp02epumo65Ju9IFdD96ScRiCc3COITc2q
YMAXIR+x1DuoN3a7RuKyghY9tCXUKkeEM7igMMo+s/BGuYa/lo4N9foNgH5KfY/8oHRPQ1wi6k3n
FCTJK9BPuEjqwil0mAXpTUuxBnDJnZfVc2+EAATsprsfIStwkYe+RgTl9z4wSW8rFNuSy/wzXmPx
ioZke+4QzfuLaBqP1SoxQL+xs3n7UPZ0qUZuztEUKOUZFF2jZb6QW2IXMcNkv4e6Xz9jF8UaElp8
SjhrJRZzXZIaxAEC9K/mchf3WY7zx+RnPGGJazaZa+rjA0b1eqUJ1aXrXcRlzeh29z2XGKLAr1HG
u3b0XcZ7NG9rvRNoMWhsW43DoeVPuaYw186J6F8zdCRYoOESDR/fyB6Wafojt3F91C+tOTbjecP4
r5mSCvfHKZUYaZRv14ySV1G7DExGksZOhpbw1iw13lK0vaS3Ygfbqh4YQTycapgn8Dn6L0ZvC1zP
H/M5pkyyJdte3V2T/tlLbLPZ3btV++yPoaxpg3lQ6HU4qz6mzCSLRZnT17ri01CWVMhQF7DJ6ODd
ix/dZuZve6LLZGATiXQmuGCfh9PQIlGXrEvHzXxxl60HU9ovXanHD5bXRRfTzFrTa9ipQZC3wS39
n73+PMO1rv/PGhMvCV4CztJm95izChAxSpX/9yhylclXezxNIynWEaAEyJEe1O3nQ/Vw6piWGZET
UPNKYAlrE4qu+1N50S+GXp/pbNvzm5sRqvn2Kt2Kk+xu0wMlLTJNOFH+InSiaEyuFhwRgMvEH7/U
9NJtqr6acVQwEYRQjBKwfZzzzsnKELDYVnH8IjheKqS27ARLOOeobBvk1lnAX9tBhjbfuMPRT+z2
kneNtkyJ+59WriTzcEZQzcZ6TLXD5p4U3QBsEgDmtFyWgvzuHc9XmFQ/+qR5ozBjzH4wBubwpbQV
8SDNXFIqCj7Vhq4E8pdO+qXQ2YcR39xyM8jg7BLZvHl9+wawkRmXJ10HnVv0pYRH8W42I5xGPACq
w0ueQ/dwupx3XEo2Vm1Ld4q8MmKV7svQRMnYSXgs7T5Ij/vnYp3YSXoin/7Xpdme7DZ1wYG/6aqy
7J0hFdXcHf+rUlFR0MNbyqMC5VV54GL23uNygx+rqmmeWTIshlmyBLoXNFjrCimCx3iP7PnimcPg
Qy4Nup4pJTjzr6rDWoFQKbqlIbnbLLRqjtN9jGw5pKp0tnMvGPn4nM6+27lznLG95cmhgXDYZFaL
KGIxJA9/L6LmbQUkxzLgjsNvKxGBsEDthMFSUCOsE+sKihKsEYDX+4ocqOS8GpJaXnWKWfQ+ctfV
P/ix3ZKzYUKCvLypgFmG1S1D/03Rb6qkkLffdCTtRq1K0yH88dNaIH/wX3wKk1ZM8Un75VF1T9uV
04wnfx3YP0FaXO2L2NZrQXsKda9uYztE+beooDOANjiux6Uby2hzx3PsuxvW9IrVo+tN7L1ig/Px
O7OM9wuRnCoeK2O1m8aWhZutoXutaBG4XTqivjYyaTOoGIhQ6672NY0Fo8qqzVkvut4Hg734Acqs
sHY4flZw3LU2vCnD96oaa2GfecCNlacHrjzDNVlh2tMWK1iox7o1uA+xct07qjExbSS3UUr7TmRZ
Dyx5Gx4Z5mApHO5xcbfo6jHUF3jrrtmIEYjU7Z5rDDIYGvZDA3vWB+YMa/neJdtmw3prWW57nCoz
r6KI8m8papsMxruSjzNhNtDzmba1H5q9Lvi2X0KEevQPBxxiKYaPNj3EaEDj+R/cfsJ7ZvaYOXbn
hv+ouHyNgJqFaByv+ErO9jpKp0vMKKsBjvVnYSivpEKtLB3YuLFTgdxCBKlyWEfYwkzWP6e5btHv
P//UKIJz5h95phcDea4Z8hb6hrwv6ycT4oVfP60rC9YHgkG8zCYQq+EyHO5gJatIF+PkdRmEFMqQ
Z1Pr5SQWM6lkBx76eEAz2my7TMuf7ybiNshjCR7tEa2jpdBImEvtNMDy0GZQaRkjdLasS3MkwBQZ
Op4VKTVbjZn9rG6eMekoP5gsnssQqHOlOoP9t5mqujdBAhYBaXeejz5Pf4BsXe288+BAmrLjiQDy
1hFPH7P0JQKzc+bPJWMeizVkQsvewOwY2RKSoO2/BFYNHEhsGD3s8QB2buCHjE4c09D3hFbgijh1
6ZMILqOnZ0ulLCxCzhPWe40HuufNb+gAVgNT80VWfbnvafmcYgENFOr6CeDDOne9PysehsGGVmqK
SzST2D/bIp8m6mJCJC7OwevfC96Lmg5vPa3MgvJXYi/2AWcwlqUBNc6aw/LxXdErdeBvr4Cqp4St
TrkXJfasvxtRoDFCkWpbLuYuw9vYO1p6Z036A6UewM5YRYiZd83p/2TP92mbdYpQV03VPt4ucMML
ZUSoqSRzidjnYC8GJKzXW7aYHHYTd8llgSjG9BSa2YjtydyW8ehyFfgvIWqna1gJ5MTq9kn+YjGU
u6VkgTI6s3skASiPnMn5N1DXW1Wp90pKkA0AYN0AZB7f9khQCfHy31Wd/tZou97X7R07QTPmwLyf
m6jZ2LrLidYRd+REcUqujJSFjGhetoUldKn7cmNCPrU8hrAkMTFNesasDke73iI3EPXxw4hlAato
NJa76wNen5uzjl3dViaCIZqV8jwwfqsFcmkAEm8jHv7ho4K03sM9j1eFFWpKKiJeQkLsEKuKel36
J1dK6+Wcm7oRuhIE+J+avJ7e2kng4xml48PEW1l1M1gL3TTTz3TtqjDjjfuMFny5pCbsJO3uJLCD
Rm8xJFpbgMEW9D3ZFgb/9q6Lpd/AoLWknz0DUbscqFkpjvj+cjOMknOarvVtjlyyvJgze9KX6TtN
5f8G/LVgWVNTx8LROm6qbqPSduDNAqacoC4c41m5RojXniMWWM4YEI/2LIE0jSBzm6EExNbE9Ybs
HRftcvvR4s46yQh60SFYiPnT0b5mzNfn5GusauTRG8OAss4bdbcSP6jOAEvlmHusUR6D7BP/3rFG
WbwHjNr6sSWEmyxcFpkreX2F5GqzZ6s7qyINsARSezSU4DC2BpwXnu+iEprF6pdum6f6TOCa7Ovn
DrKVONZ6Nc9mrHRl8XxRJONNWQ3VL83hwmUbxAIwG3cikIqkM3ewUXYYfMJEN1S1JE+pkPK0pptC
n3zrncE5Lt8oBwbJm4BkDviPmuDSkdestv5rAU9P/eCHUoh7YC+UZkC8P1tuFuUxY2r4gbEJA3cS
F1cq/17/hXIV00UG0oS9UO1R+u6ELPw5y0GJJpshvQL3WQmu0ySly1U320aLbw+FfrGXfjeXmWC+
ALTw0IgaLDwI3gk63uPW+gn6C6i4fe8PGHQxfzXTOvkqF5c/IgGe/Gsg4zUlTo6Lzf+pySJX2Y/2
ggQdR1pWY0lIZOSmoO5xI2FifkN6lk59fUMyMHYvNPpdlqVXBE9IdhwHtxkOpQbus89YqpZXuXF7
WniFSE/nQuAJb9GM9P+8RLDwOxsTSSYy17YL6ejaLFt6OvEnK/uPCRT9cjycVtPYPMpT7elLH8Kv
rY1URZ4rsvzIQRje5usnnd41GBH4L94BVuww8DymQczU3X0zdo5Cfv1OTE+HRTFx3kyKEtfCloYN
013b2DyOnRDASPIx1NCHliZCurpp/H0cs99sgMm4uYr1qtfAoj4xE80hGtdiZh10G6uTDVj5dW0a
2QhAaSoXSbVasoj9morT9Wv2YixlNQ6OzaX7Yqt9bpfhTDdodIH8Erg1d4OQjZEqbhakKmGDzUdi
z0LLm5Bfu4drYl9XCE8mttOBQ0EqWA3kc6y8QgaPIcYbctJvFiRRNcusUTUBegUAcGRfbR12VxLV
LhAVI/ypB2sagiAuuGZhATYlqcQGrc1PNGzR+V7up0DakDNl7VrZw6O355ahUbWzAXmM+dOom9SX
levE+HsAwhpq1iQrtQS8c3biZzmDuJPDQtsWjble1vdFxa4SlAn2qAOaR6OEx9z/rnw+zWkJ/Fby
R90hWmjP0Gz6RXgzd5LLgbwuhdxfxFe9kQ3+r3Y/FUBll/zCFgzs0EgNuVvZPfmciXxnYx5GA4XW
ioer98aWr0dBNR31IJxKjWzPD9loZYfFTDGUtL5nxgPj+rCWtEm4+QShlYaFf5NeR2v3DtgWFi0M
2K50c9f8vFkZc6rBQAYDh7RXOx3nU3sBYNi+zQQLTaQWZsjbcN00+VsEtYyVZC2b+CqXuSq2H2Om
KJLSc+UM8M9GkqYvR20GeeJA+qNpbCFDH74li8/Cu7nX5VD4TkHofkcsipWVRlFVLcHV63+O7Y2r
xXq+zsSWBaZL96pvco3ztVkqjXxQrmEOnH5a3eiP4Pw+knYl+Vi1Wf0RHTAjEMs0TWnEIAaVvwkn
dEfb8BbReKRib+ZW5cTQjuxeo/n3qLcusg7QLRfF//BEKPvl81HKWiysHHMlwLguahaD9hQnzoZl
dFlAN8ZTY+kXgo69ASYXKa0aXHRUabXXh6ybZIIhN1jsgVSiDDogvOChlPmtv3x2g7Z30cMBEip3
8PnDhglN7ZbVpXZL0q9jbt+QU7DrMyRu2RAjPHZ2JOltIOwVCY+Iky9+TTnw96N6vq16SLClUvZQ
BTPP6qpspV6egPu9ozzJPbsTwjWTeqOkPoe+mG7j8fXECHGy7l9JiJvS4A2fvUw2Ty8XxXwW8KqW
pOn/g4sGGGeUXlsXFtY+mYk0Y4igWcUbha47t+FZ1o1O4O3n4ZB8VcAtmTDOYp36BQ5dJJMxHoz0
H6PQW7q/Hu+49TMRgvfgWhqFr4HNWR3hCpSn82TpqnGGShhJask6lx9CkCVVup4VujAL9KeSbgZf
udSXXqgmGeAr5y2qr7luQZN9wyq1/RAlmrFY1x3ht90Sg2RdjlrRYoODKU0U7Ug8roqDAu8O3REm
KrRsFJJe4VEh7r2+6G+pi7bnuufNT8XXI6D5wdYPJQEz0qOV1vwY+ICgCeyiV3nUvCkSeaViee+7
tBH9wwcFdsU0JIt2GpK4gw+r5bm7mzVq9e+Ad1N1DLfZpfroioKB5h6vjxjdEgjIQN3seYrP6m8g
UvL9Ybo8J9P/tfXbMIc/pURg+nSolSuk63uS1labNu3ujocgKGHP+Hb45cZjB6hsrJooiuCclet3
3l+2ziXNLMxtKN7HndBGJ1pI3bEPtAqJOUELII3PnmNK4DrJkCpQ99xMdTgbZbGapkij+M/78oF1
0gRBExgjkTFlqh6+6TDw2qS0bNnTulAPehJqBsYaalCk59CtZ/HSAuU2h0t9SqheqAtIalqmpfAE
m4iA+IiAmwCNY/Gvp5TYbfqHADvs+rwKqZoKQoZ5uTGLhO/rVqsIfr+tCQhcbkW7HKErxpu8Nyfu
IdgtysXl2R4ZJAuXWPzxcc7xeThT7pzVyR3sRpAkt3+MZzhv6VqF4EiC4h00rKfpQIGe87bmy8Oy
MCKOd3VQeA/fuSnyk5Yi8tdIcQMuK/zkhdY9DcnplofKn/uvtq+pPklTP/h3JiCNOiSvskGtyF22
2NOMxyVdk08+1PXGv6BVh8kv8yvkQfMBWVrOGXkbRSnVVg9rjSCav17YRVfihiU+qXVgKaoRhTm3
pa87OmP22hDDcZiD+f1etJN9ijI3/YzGCxxDZpgZ0Zx2T4ozFrsswZyO63LieUGyBmP+Sl4T+2nS
VjNoEpMGPgNrS5nHErVpPQsv8X6i8h5vTmhM3Boqo/iY3fsFj5BEapxB9/nej8xY75SCAteRawsy
Mf17jvzTTK+duXSR6cuUkKepV4Ex9FVofCvC25ZWXhwRgAqWBZ60GpKgwFoMS2SCf7PIyXyaIuCh
BzFMyKYJrRhRW6sUj3nxptcxtRQrNSPUjsZVjWzpHyK9PIvQYX5dxvA1JsFsb45XL+LsjjHRZlsz
SxvmrmQM1utT7w70NbxUslFGl5EMqSlmjFd9PQXDQuPqKG2+nHoNLQZa/4catm1N7j/9k3JDBXIE
U4QDwW5SFJGc/ePSbmWyLrrH8ScBOfA++39ucGhz7GPug2Ea/oOkYP9/kdSQfReDm5qJN60eOhnu
76y+OejxijxNpARXoPeLaNCTfmZ702XA/bbtuzDzRmBzzIbET2wyD4JQRmmg2tBjnURWr+h+jOll
70GZuZs6D/W6F0CxlPH4AAS8rO6M7wzVW8bnfWR3XlbK2TvXWTjXbxM8DhJ/OuUUjdk5ADJ45OO7
+rXX1IlaN9LFXG+ut5JjAKCcSN6esTkG9VWfluXHWXi0EimM71U0Mfyn/x9hjoS4qllFypn4oowL
jW7ppNJKbyqPEVFrt49iyviPQp9ml4fvUXQh7j+5FKDs/RsX3M7okey5m6T/UTAx4WL9y/DFALIM
yFHWaI6/IPyYM0NxQVtnKaa5RPMMuYtMLLMaHuWYsRt1FtQAejzrzVjkM8+wPn+bdCTYNz3M7Es7
vKQ9DvhGPeBgk1t6RPJjSCpoobWnpPeULXMqAzeGwBAt+DCQ7EoZCU03cPKdS+NjBO9GpHKuRnSA
4NGR3uIt6RwrgHL30GhJ3G12z6Tfty+z9qTUrkDQhaiUQoo8lagYFvSlqv3wSMdkLk5qPtN+BGEl
FllyeLJawyudDn7IfiFpjZAgaEdtvQtRxogApULUhfsJL7FlpGEJ9qVJRCf8sCmZJFu83QrflQZ0
kYFUzqs/SfBjibtx+PYPqdoQdXXfHzi/TbQQfbMJN/Gk2DAbgypr5SH3Ztfeah8IvR5RRW3dSThl
eRoak6AvUgfaVAVXCEyyuljUe7jaGZkWFkCCqyKa+JC0v/nRgStjJWrJUGYHFZ0oribxeYA4c569
LJBjZ0wtEIVCrb/2Ure4YHp5z5Z5nHCIS7qV3PtA5VWEZuG5iZrdTKqenzw71t4YM/uOVNYxfrXK
OLdN4ZYDhNoB0YjFeH0FcOp9m7MJcJ6jocj01Z1+7FboZgPENXE1O9Ix1RFebv/GeHzZ3lSFbfJ0
iVsFluAYL8zdP21FeqtpbKzTeni4O/uvFj8CEC8qsDgJVD8SZWQrLqA/xkSIu0KBkl63mwO31oW0
44PmvY3y4Iq67cciBlDXByXAKqOK2saAmpG7/UHBHNzzIf2dTFwEhKyEKWjdSaDKLeMFmqJdtGEp
WBRJHBHATu+fJLdAcV08l4u6LilOWlDnli0lSJFKeRZI9LhwpyJeOCpYCI5u/luvD8qacGm8wEoZ
GXjrbUS3NREoxTYvPEtbPpbyflky6n77aGI6UQdKFRAccdCTwCBHRj3TfdyxV4axpbEhZREob6RU
ylNVSxwr6lkqXZ9ALwniBr5ISDUIIKhlSoIYy/p4EJBHCKbyUXSFd0guWtfnHk69OVQYqL9bFHzg
1xYOqLkUGIvEOmt4jof4nyG63iK+OxGF7DRjmMiyTU9F4NBn5PXalZTdkJVi+Mo5rHQ46X0HZmmg
49sS48AhB0ouIyYbIUvsgNLpK221PzOR9umFPyO+ZGyJf+J/hEqhtEy2QwCv3RADCb4kz+eRb67e
c6zTow7qtVHHkLi4pPC6FcOX1K5klNSG8taRATZ6y8R8bXVwJxM0g9P01KT96KG2+Brw0H0cIvxX
2xBYEZl0I8bYFduWPsQX9s1svQbyvPBwhXGu8Wy3KM+t+zjxIwpkoAjtvzYDZ0O6QNGblxWyAxEU
c18T12gNmd6MLPkS7uzwefCIsNi9XnddFPkL+e2wofQoceRstg01FngtStfG/+tM86s69SF/5+XR
1KRN8s1EYeAwvAFXkVLwHE/doRvLJtwKuUxs1KhTJj4kNkwrpa1dPvVY889YBMjJ8f59vRInXUWc
gQWXMdEnjFK8UcXoo6jfUAvO+QJbLdernfvzwUVc8LO4qxD3ckbz6hD79G2Nu6RIGGWpq111vTFl
m3gtvxBTQQ5SpiE/w2KPiSstuVBPfePZDy80L1NmBard8FWO0kntj4P/qGHoTMPk7r5L1ERY1BLQ
beUo9NOorus+FrG2UAHBkEVR+ws4um9VnW19p89jAobNn/THAwsQFPT9wCIJ/ACZ4nbo8KF9G+YP
7/8ZYD2u7TZwIqiT2DiAjGU4tWpI39EyOmRJL3BnX8y0eS0vB4yUzvVFxsQE/HEEXE3zP+cYmqwg
vQf91wCPB05h+bE3LQ2Cc6GEvdrq/2iLBj10nWuhT/b5dX40rtPbpbqqD9Hp3XSHwJ8VeddRLwmc
4N5GdxRplBrCWlWVAkNh09gY2tQql8V513uQ7QgkclDT+9ZLiyg1kxsl6T0I3JqD1RrXdqZmQKdY
m9C5aNPv955PcQjnRWP9hkZQdE1Cf5DHPAXcF3z6ucy2QUUoP8M5M0RKPssH2cn4GK+GA44OOjcH
mAETxuKWIcYq5eedWYjS5pnCVC7TSux03Z9ulk4dBvkF5z3mEGgaKEJW9uaIiBvrzr8tAmuDrbGw
+jvQG91aGnhFWzEZsSwriEG8UdIwbPomqpNoXVTp9gftFZSE7vKql/tLnvCvm3tpdHKl37FFN/5m
XR4FTmpi5wiNvwVEfJ0YCcVn5qKWumbOrbBzzMvQGX3ZGQKPfeF5MQnO4KkzQ24UoDI6005oMK76
tcN+ydpMnKHOpscft7L21MSMi4F8Q88vWd06bEq0qRjcK3G461tnq96+8FN5/xsxhUI8Q7ahSREE
5neRQesBCEUzkqCQjW8U4SV3iyo/CIHYfmY59bIBT0HIhsqVLqrqXS1GZjvUwPWjtbukJcToLV5W
EgIBZLIe7d22Qwok5sOxRzVBDZuSOFKjslKEem2SWnBjzpfIhZAbOrdd+f71xyJH45l3+gfoT8yV
yYPL865SFlwV/Ntj8ALTDZaZvE/edPFNL0tSV+zQk2egHv/3pWmSqKwVuKtGDubZ8WcsmHppvdyV
kvPB+WHZ4wCTi27Kg/rNA9E1UJ79uAw4uJ4SXIudwBP+6rtLxtT2yFuvPKRKl7g9SUuRFqznytq5
yhiOaDq98+78VPVld5GESAEWtwpjrqSjOzqqd+nXnugeKkhdCPkAZWE8eGxLq+gr0r2+luCrSAJp
YiVQbyp9iSNxvXqsxmjdydHU7y1f8+3HqKjoyR2NdCICUNuO0os1r76qW9ErdQq2Kh4VxFhBrrh6
lavlaCuzuMq0N/3Q64CrlbEC/pXUHjfzvmY49uyP84UFig9DkbCCmQZUMe1BOqsDG96lgwymipOe
JcZ38+dsLAaCBui+74E2DlYY5yFkzqQqXF6qW9lvsDlh9quplqoZuAdIe/KdubgjNjcYNrsDKrvY
SHTO7lNXSbkHlLTF3PgW17cgavmZJG2MyVarWwcgbLVMQqEA7LFzvFj+wVktujJlUuToeGiXO453
Re34Q7efVa3JUXS0GNPjmuTczH3gLSPgf6OfB0WSNyzf/AfBn6Z0uo0zNITl1cEV7uJXR2PqgQaa
ydrMNeaKv5uOKPYvsYDK6UZifP6XUrlsNIjs3rJh6bEDtnw4bKMyJmvR+zWql+ZCt/VCXyHxRFQM
eBaDgJjNZ4upVU/WCbQeJrQsvGv4KqJB3azRGeNtidnQfh+ZLDJF544uvqkdsrjK5GEyx4jAPqtn
6tNNRl9+NLDHar42nrL7MuAoRI0ZYDSd6nkxhNLrIOf1TH7wM7Ehuawta+Os+e8twVzVOC4QXNGJ
Rez5GMjO2ANzeuZu6PdfU14gXCbGVM+zSM76Z64Q3lWD5tSEstlUGKX0ivxfcIYHAnqH7VaeMGa5
ldJ3HDaEjXLV8XEIJU9evg/7OCRoI4Oyq1UDZsu8rze3c/jOH4VvTP/I1bTTDd6PAmAZVpnl8S1T
w/+Lub9zjGbvA0hpJ/bJzdhcTqa0rFV6HSLunW7JLQRHM3CJ8hgPAWEM3MfcIPUefZO26kyN85/h
dXRLWrCll7FUg9epknC6iPZPE042jcJg1AfSD/GDZN6Sp0setTm58TuXxTUui/eAJ8kCW27eARBs
ljDZJcTbeFqdqgIMe3Zh/L1J2vmk+h96xMaXPZmywb8et/K2eihSPT6lzVHIP4j/EoSsZQhGEqnd
LctQA9XyRphiirUszA8KM9oY4cz3Le869oJM5O6aUbqqnXwMJi7mRZFrNZHbQPQg6NNIKAWbPsbk
gD7nT3j02VjZhBQS88RPQoMr1WEx/Xybm+ATt6C0kKoy5f3q64nJa3fF0mq8bpILp4nGkrAJjSc1
cu3uof0Uzf5TXRLLSeuUbFIhwlUH2CldspqLDxyqaiLDB+q+BvR5FwnYZH5n6vUzdhkTo+gW1Pbs
iTeNWDMbpsv4z5oiTU+9VPKewmdDB4VcyV3dal9LEMQAbEOWQuF8tnVGeH0/Q7c3247RWC3BwNxr
RFc5/xRjEkJ+lR9fJX5Vahoa1TLlKCQOLEBA3dtGR6vXA8NsrN3k/U9cjaKaP3cfEbdMRikcQk26
SJr8thFLahi3cfn1FT+SNeLueU8rEZupKJNebCcnqU3Zvzwko8SDM+1IN/1dJTTrhKm6W0Q1yFiI
GHt1ru6y7JXyAU+Y3Vb9xupuzinpkHQ/UkV+jLjG4DxfRGGz1RWENLeZBeoU51W9PiLAOLBTdfKW
oCyBL1pYBeyoBvvDXBbnShA8ub06lo5JdIEAGdHN+sLXQ+LsnHyGAvKTk0OzPx7bgewEC7oZs08d
rus1JiG0ZKTyRWJeDT40T9rlWGc0g6C0o04dkEHNJJJ3YXfsGpffRL7OoeMAjdt7BmG+0Z65ZUNG
vlBPT77+UDC4Fm1HAd4qEfgDMlbaRCr/HBluDgmJqZC+Jt58mjWpUV+jKf01zpKbOe96po9Rpdm8
+s5/YIsSQTL903+6f6UkvjtCAjT7Esxnnqq62W1Ux8SFJwWZOZEWt06zMOVF8OKDqoE6A90fW8G4
8Ci25uBlBqxjGmDCsLObp70W5sN8FvWzDpDUms8QOsgEO+TksU+YFlXIpK7uXM0PJX+ctBBUrUNQ
iPtAQb14EGgwOintbhaqD5PspN0vI/PC3BHIUu25Gu2tWxkqqpx4cLBb6CC5dBgSdPNeHz5VyudW
1YVXblSUOwoZ3LIi+PBivkZqv3E2yLlsmSKFOoWmib5NlIyxZPKa6ni/ahVRVQMxuC738FlGUHuP
Ks2wbCDJuAIzTDkJ8s2ytIJTSXGYoFfQdVi0sYiTVXvgxWdyG7BYe6n7YnC2OcYNk8rqNow6ObCP
ZH3hvfzEwT8L2igYKBdOBs/i05os2dVxceu4fPYh30KoqR36GuaBn1pZ8ezWy2F1x7RupfjT2dUt
jfFSXfYMsfmY43vzFs8Oe6vE307E8zswHYkYAzh3rjr221OYKrJu5zHmp0MkzDckybLd+gfgmbOj
vdAA5MNrJ6PYhSBdbPAgu3diF8gikWhfpUrfxzY7/0yfUZRtqjR9V/70IUU6ZfIZ7bny+8NyDBCp
2iI4ESrQCa3PA4JzjlG/pTglfcvv5N8BOzCptx15s7fXGitn9ivdxZrhOZo+Biw/+sbKQ8IF//54
cbLNEW2ow9FldBcsmZaI558xyDSD2JUKPxKdDdDfNUm24DlMSWZWxTCXAVagOiEdYkS30yxejxd8
qAMmRzbJarWzur9AhB6FTJ2n13i4OIeH3CBxrYO7wJl1yEz40YOgPzMk/ZyMmUoO5g18FNzIp0Wm
wMFKEqzvRCqh2UckqhTkg6o2D1KBZivqpkhD7tuvmJ3NbZCh0myAXEPj9tizBLJuz6xEvbggoz/M
Cu4rLUoPKNkdaY0wO+SuGeY/glZclctAPYvAkcMaDQpI04qlWVjsDz8PsggdHRypJTJ7RWEu7MDv
d58CUbI+LFuVcZl0L/0Aa90SBAdRniXMRK0cDClaQgUBzqVQrVqdgQj5lyczPw45r8tivjFbHXb0
5ju5TJa7lUbmH8o78MJuHMVFKuq0hDn+shZSnE50oP/pDecxAhlTVWKKIGA7qcDdESD6q8+9bahI
sT150VIjoXwM3TxyaslPiN6Z0oLnwuyjsGsUQnsbxCEH0Wg05/2+8YYjdc14tcRv8UJTD569LK3h
EHU39xxbp0D+7d1HGfszg+xGHg09fGcnm7x9JjXACVtswQ5LvUgUFGTjDNSRigxAWYM9VrKx8LLJ
K9z9Os/2X9xc+KELlOce4dMDwL49H4YUj5VrmY4oUiFlMe+L2l2uawE/EOPESa0rDTTi7tYATPp3
ncSWkDNIfkbFbFiSzLX6cHBNtGv1k1tEZWI66c3kQV1LesephP5j89WOfQ1OpIrtn/mPxMxPUUap
DcjJ+mXuLDOfvl/xFZk/Lvb+G/wYc4aRtPRvxIZb+DORDx0byPt0MqDlZOJ5d9kYalr7FqWn77KG
2gEmZS3qX8bhHKwMtjRgMbVZZbdkIIw/kYB5rMHiHv/5/Oa2qrS/43CgYgpS3G5zf7iWfeHkp7z7
KXRJtjgLdaXHW13/Y8x5WucoQgWP1VL2BzNrStQc3pL2GOgLBJyAYjpLPVqcVDxLsp8iQXSxvBzp
0m5Vv9H6pUypocuSFVqEyxTc52jXJpcp84KeHHRNmvTrSqsJaYMEG6+STKg4wE6KZPneHEVodPlq
lwZbjtXlxq7DzkpNu+4j4Y4t6yFF87MSTCk4fWwpClqsfQYyCf9BUb2i+IjS9mzs5IMCeJsOqwK3
f/fBc5kO9I9MrzIKAlzbgD65WdHyktATBvsoIgN6lL42S6WsdpTuP9jL/ThRHMebhkbpJFSMX6OZ
ez22DPGyWXnu/V3EfIxlxIIv7pSV31TI/7Py65rLqPG5t6Zhpzt5aRKjV9W0ZO78W8eR3N+WFvwx
TTLAqOZcbFf04XWstLmNjC/2hG4OBGMgqO8YlGl7HeZ67JHwUjnDYuxjf0t1zYIYMeYkgY6JHJrl
Rn/821CF/IaOmd0zOH6htMlMyVbwkVZChgnj6uWQ1artTPIiDa/oAUWWcsDgg3tGtNl9Qe8Zob6i
xwJTb2SYT0i25goJIVwyWMLuKxOJ7mbqCgmK1Bb6urSUM3lb/CYksSQ2nh+UDkS90P/eAW0LARn5
YAXsFARf1r1szEJYSK0eF6BWZ6AYNM4kxpQP0ulUODtgoRWudVZW0rwo9KccIr2WOcLxxT0HLjcW
HGYq24hv420GfwPmmRqCqUkxai8je8IGHIjEwbhzsYNn6IHtSmQQdOh3Hzc572sAGV9HvEOx8Sta
DtGcj3YC77F+tp+H2bbiVO32RAvRQ48C4Z96c6gM/TM3SFlC8ymVWNckkXx5gDXvb7LYZE1L25Xu
AK3DF/BVmAkytr/R4MvmXugf9zFnVY2IQiBTvZb13ypLd4WHDRVySk3cToPSPPBg/XjA5g/AyBlI
wdk7hIXUPYuXZS/X4lLg5ep0B7m74zzTxGVQCk84O/1QYtDeTAzXG68N2FbkaoGtdohvSq36OL7b
YyZaMqGCFrzgp2TgpBG3Qf9i4dC7yXB601dQlXxRp6Ju0ER/q9oL6/cebJuO0K19gMsACdWq02rN
Ckgf+KZU4tSnUBzqfsM/U0a4JFKn1ui79jv+ADSKS7ZBcQCU+AV7Mmei8++7hWlzAJJsR4WVzzM+
7RUREBFQFC4GQqGLcnguasxEprBErKUKM5y+mZ2qYnG67eE+CzxrF+ih/xuQuOIxKxIqajdKCdP5
iRN4EcQdNx+WSTY/44dsk3bIamgUv8QdPU4gUJwDyCD6+DSoWj8dQ8c6YsGG5XgAV2vm8oWSMxjn
yUevW+wViwi35SA1eL8zLC15ywL90LwnnSvcm2g0Iniasfelm8gqT5ONCBRxT50YlV5j/K1yPISu
EB4We06dSr9y/HEQ+2qF7yOVbqEDvrpCeAjAcVRXtoZ+41BEFRKZuoa98w77+iDVEjoIR1dJl0Fr
yI8gN35EQX6/DAROSFBtJZabGCJC0s7ynpsyVN2D6V3KlR8wgKkwUoWv+brq4yO/Wvg5ARIiLxU8
HIuhbv2xatS1GgW7P8ZSOHJtBrzqP9mPQYRl2vfUyv6MwOzHOQbSYV9QNdoYSDIT4ZrIKw3qdQQi
vfCZaQ8GmdLwJsbJM8ZO9LX+5zYa9Ry3fxjcE2I3ZlvlGbrBp6+LGYKxI/adHn4GMj2h414CaSR4
Hgy1QqfgzjiBAebt9ISH+Hm0qpK4IvLLU76sSdZ5L00csFN0QWOnNKIDiHpqujUcWbJpqu0XRTma
bjyPBAskuxXdVVZYtNtWXdSpk6KI8cKkByxgS5LttKwf3wQU2FSQpfLzKqo4kGra3pNI2FVoeeqL
xZmFbgNiuyx73dhyGD8Hjjwl3E5Eb88uF2wCwEJbUOLeWqMCiq6GipwdqUljPd0rPruKgDIVLD3N
+Epn1hw1H+Fi5adz3NcWYDLCFAe7EvmauMsBGxwAlI1RWR25eU87O668eLhrExaOJSIA18lD/GTJ
uAuXDg/pOeIYGNpUb3euZYZtiZD+DjAsy0gcFLV7B+NdeChg/Jjky8M8cnIR9qjpdMWCHmynGfz6
k7QpVOdP5m0V34LpnrkVLCTaR2kncqOb7GXkvltxq+uSDKRgKyR/zKa1k9taq+oZC4VMGXhU5dWY
vnaFx18igzXE6FKvsqGQ7S3BMZMR09/Ui/j0CDXsZU3fKPUpyvJS/gHhTa8jdkV9PASGJRNzkMdH
2y+3ihve7nvG2Wz0yyRPyDvo5dMzGa2bm4ZDG7DpYxWpNRBz5McqM6clbNxmnKvZRciZWUjrPIGs
nmnZ5oGyHKdd2UWjCE6S3fAMAM9sZHfCBDhb6fFOtpCUl7rOxBRNZiKvE4g0YqrHszwmb7FpsyHB
XzrtCBiMWmr+BayKgVSnRKdAo/oqM7JWKGDhv2swBUppxODNAsxERcEx++lmYw/gFutXnc9wnB+W
LCH1yC7qp4Bq3Kj5naDzaQoXgkr6mfW6oGQ9/fgbG8kYGPO6DP1qQsftmCpWbiQydKwMPA/Cn4ie
Pf1zQHjMGSyV7aIJmOd8VtontWXhyzsJnr916G9nrxX0Me+k6pO4cdjF1qO9wm8Dos1m+HAFggvP
9SD8DuH9WW1bVy2fKDWLcTb/vV44xDdG2x4ETbQchfn96HIFb1k5ezr4aOTXHvfw/HTVnvhBtBkh
3NL6GsKc/d4NGNfHT9TdepOfVwLQEw3S2CeH7mxOo5537f1YoWvwWgqXfj+1aGnOM0Ye462rDFSi
SfMyieFlUjKhBvPM+39zZdTtZy8fkkBpVBSMaILTJ51vR5B7vzJ1p/0HQv7nopNETdvtYMyiAlUV
635sGJ9T9dgsJfOja4hiAOJHIEm+7dW8kOsu26+Trl2vHAFQwhhqt3VbuQmgUvPDpYM9sBSdRWwF
JnHKvCQaDW59LERekW2ah8oBTEuApKbg6COVkvDMk4SmccmZC8C13f6AclyK8PFDEMetEhiiq00J
nFjGk+jnd51fyB75QkV82c+mzV9fagFPkEYqvdRjIjPrAHdyUjIzDqalcsVQkm5KBgKb7gvpJIcG
Qv3zP9as+UCFm/JbiNYaGiQPxckXc5siE009npnjMfmELOpbPL5V2Tx9s0V6SKzUhSUJsjpY9KV+
x0QYmYJ8ItX6elV+r6UECrZ9+ppd2h/xQ73mnlDuPZoEKDfCXcuhWcdDRhHrdgaUev9zz5qw7x3y
SL5c4184oBdQVLtqIvgIdwf9+mpUcqd/tCm7EtC33TTTS/NXkN2eUr+fBBWxO1gaWCkhXTh/kSvB
gFBt1ZaAkXO6EDT4oEm8VkWiYtI86RVAecvfT6GzJQn6PU6/+HoXGsbJtsckoGnRdHJITnXutsjw
KWNKEfesHvk8YW3QBScWzINoeDfWAMzrKNDIvOxyI1+D8/xufAOqynlTOBTkEeWehQ2zIDop6wRG
Rh2gB3Zz83Eeb2Rx0xHB5rebM465xlA9wHNow264vPdwjZBZN95DnUo+ES7yz3Ay54OmMDossDH0
yZm986IYoWrNYgQXTdrMOoyUSP2TQ1yLor6djkotxbaq9fdypfJEpuv9tXCavwtGo3y5d/RMm91C
8zVoYCNK9uuTe/hzYgjCFwhWjCam9QlBXXNVbYmtEDPmsabztlyY65JnROrdv8kOkwiL2ZTw1ugw
6VPPHBd02kXbOjQpwRK6+b4rfO6e7wsEEt/ucSbf07KhxY1ngpKpO4ER9hMRK8MXgjUYAncy69P4
1w5crv9V85TgXw5mwswYH6rA/pkL/hd5t51Np0tHNxWr12MFFbtRTpuzwysSIewSa4wsSSEIi5yW
KurvjB6NePCAEyVW7vulfHXxEwczVAjXBl6ZSZloY+0IBssbqNUfhG3b0ophY5uHPVybf2U8Pdfb
HElo8fFxwYa/dh0svl51TrJzAVVwUmDKIoZDC4s7neBYvHXYjg7ktC7zsRdN5SeqjDF7yPVWWQAF
5TfgJ9zBkavF07LlsWscnYRZcBHgy7fXHNkdIXGkftuw/low0zqh4u/Ev3kchmMVvnRAS9Dxyk1O
Bb/EIvwovjC1NdZIm5jGavs/Ap3w6ZoEfzGxDxTzgMqzJmxuUlyNjjQ6vKDmIQLL3szhbHkhxpuu
OvXcd7FYolLYw0qyKSu725HferkqWXgZ4GZl4ufyxjVASFQgTJ8R5tCMDzzUaAxbfYcWqZA7YeFe
OVZbFjBim5hEcYHcpPR7AEkyK+DzimbSNPn43gP7l3joprSvu4gDQvp8tYpHX0GivgSnz/JbDE1o
qWo4IkEL37lLtOUrz5ltqpDPcwE84zZHQCgg1LvSP+lwZLOUM/pMF2t/hf0/zn+IOAtliGPiRsF8
3O+eT46sjY6VjC7OEeWtz0wDijXVLQW1aCRw8Ze3H3N0IqJBurtZeeX3K36xgQvlC2WWGqdDjnL7
Uaxkg6e7uVzI2a9gTx/5mAC8a9R0TkDYE1JbE8TQPB6wgMfX7fdVhKltvT/DcXh73x6E1yvGAs73
z+UQ9ialimu10ArU5KCCvnCRb8cCMuFJYt2IeKzOgSwu3wno/X9DtHBXEKQU6VtFGSTtSXaPdYjE
zKidnzY5Xwu1GtHttpTi8YRwIiiXbZU0L5SuFqcCVjhal//tRVr0CGDwPLXaZ2NsnAVwxOwTnxw+
+gBJ/7fsksNVXdB+776YJQ60z3J1Ord1i1kzFg3hjcg5NWqPI/uEy+//cjNhf3FQDssxLLK9drym
QdhbYllNCKivhBzta0YPCJfZaGo1cOQwJ6GTZyiNMGViwCyGW4Azlf5LKxVs1nqNroFOS3E8gF5A
MD8rokwYqMvz0hr1sWvj6D2oZeIYIx/0NHjZlACaxwN1PWC4N+8zrg79TmIQYGQp2iSlLv1+7MKH
+ewTkPcjrPeH53+N/EWuUemBshuPXo+dSew7Its3Tl8+dt+7FYC0bdw1ecDH7a3asX6IYdaCyDLL
GU92tYOinbJNTabT4GPMmhx47rEKrZ8vMAQLlj5z/YRn1vtyNQFgbeKUDBzmFa8Ym85PD/NA2EhD
CxV9/VXsgEiTqy/iobmlNBGDcPUpPs7ruyyegwX4eeAIDFr7BjjM7Q2lCmLk4r/aA4Z5COjntRY+
AM65uX4fglwY8RI0shQDaWxH72Ya1F6q2jC/y7xDlBEd3oyl6Otq3Mn+Ow/hRyiv333UALKXD0O+
HP5Ax4eujDxnjygjEXujsdMIDczbo2B1+Z/iqFAfeIPZDHkIZvtrTtxBh81ZSUsu+oBmifz622Jf
WLnlgo3sL5Og006s8LXi/GCr5zG9D6vf9wm/NFP610gzb5+arXTdAOQowealEeeBgGcIXI9bGzdm
sXoOWvTmdGAbAogB309MnR/ytdjYnhOPW1bn+F/QNnDYqu6xgR5yvJ60aSpB8WCS51+Q8i4R/zzG
8Qv48aaLtuStPhvCVbSkBbtiJRM7bgXtMK9V/oNmHMM9pBipa0WABuw1qmMqGZAlvIE3xvlQXzzd
i3CYA9FHl4AbTwRJukDm3mtGjCBp7QZe8SlMvRmVu66q303tXTXu7Wl43g0fI9O5diEDyT19niBx
mZAGYeIPgitrFt0IVoX67+sLGdEnirbHUTkjtlWum8Qebw9lMtWhlc0LuJptKSmMCcSjTSl5bPlg
t1LuUYikUxx45IfnGH5vlyTnBxGFhtD1mEYMtF1MhPDiNTvajyFwwJ7cAYUw/bnfv0LrXu2kM7uV
uafFP0sKj1IGZ9Vggao3pWMmzgwyiu/hsODDxMa9ir/y0G2si5jvtD0rI4lwxkzAG5LtilaacloZ
feM6J2zqqy6fE3+KlYAJG8t7GyROaOZU6GbC1A5qYkc4UDW34PZ5EKqkDm2PiZqzdHHe//osEmoc
BDSe8EOfSi5VVRMskoFc9nBj34+pN4MfaunjVX5vBdDHEdgDBD7bmuSL0ClkBjkM1w7qUuE/a5sx
HBuBhM1Ko47jevjRKoPjNMYck7G2giafTAV//PDiMyG3GRjL3/MfF6W9l6xHoetYD882Ived8O9k
Nd+p8k7FtoEINR8QYlP7KJNmY57O4DzUdVEsPlXXdHQX/lulRjoP2e9m+KB/AonfyBkOJHliGGwS
JKOXpOZLIrvB0l3z7Kg4yCQmBFYIKnDKzH9rzXR53ySiHtRQcR1NfoQk6fmlzk2U6FGv7gm3sIxu
A9t/eUyvaMibslr0AUDRScJczVTTja68vH3x2sT74o+P9ljjwVjnjgL22+9bYpg7ioE+NAcSOmGJ
MD+VU6iXpPkkFgZxhVGqMko5/REcaEc5IqSe+pIKHuPiDRb4v9iEOmw+xvP4nN9w6Y8hvWbYeyHK
Je4mB9mu7l1Q7VVxGzUR9iEQC0j9kGpFt5YS5SERg+K5D6RrLZCcd4cIdajw2LoQerh6xbnhugsD
cpBTdskNllNxD0oqIZX+/m8yuRatANvfCKn0jXKoyIp3F2GFiDflexWck/y80raBOtRlKlXdumlj
DMepB7rOdH4jkJ6DGXb9+ZQGU+yHbMbFTguzfOvaufucDC9We359Lnqw8k54z7J1s6meC42npm1y
zlUkIxBjYxF3kg/tYKbwhEue/9p2MyjJbIQJGf6x1ZaLFivIbqOVwiN70zyxuMYlyyq8BJ9tKpKJ
5fE6z5Vd7NP+YsxvZ+48/7qINitlfk3aitSN5VHIhM4rsZGVct1MJYH6jvlPbHe2FmrrOrjZw0ft
xHXYNltmqwMibavEi7kpL6XxlOsPLCixq+R98dalTlyhOp8UppSP37XcY1k77oJbDTZkK7AJPz5p
dMkOPfIr7Hhe+zhkNVrZM01KxfRRzHidbaJ42fk468JPQa7ys3JGIjhnHVgEKFjRPPAAumopniC5
ZSw3gMyFtfRR8cvTOVFMTxRhVpkx/YtGrEk90vKQRGt3sLKbG3YDM4HLL/AznSTI/FQxLpz85iuI
Ka4gycN6eX1nzr7umS9FM86RdMqt0hKRjFCr1M3utngE5E6q97qyXLFGXADk4AYrX5fJhxp9dB3E
kk6QRU/p675PNgJN1AO+AatqZS+9mPL7/Cew4pyIsxrrZnzxN7hnNDI9XzokA7GdLyvnI7JB+0+o
nZPbtXI0BBhPppvZGnouIBjJMv/XQL1mjnat+1tjNxl8jPlGEHtvZbhWxTrVcLIR5SjIiRGdF1Rm
GjC0Wu369TD20RYmqbSHDDSU7O4p005uSDc157ojIkBV7+4uaWL67FrlXTYpKRGXM+R1nVfxg/EH
eV0r8up6Pv9qluwmn0vpTqzdv/n1EockL+1BDH0S//Ru06HMP+TCHn68N2yMI90z3TC8JGSjuO9Y
K1A3Rqe0MaH7n1yBBYJS+UAkWAtfz4ThbWaFDf29ISt8Iu0C7ZIBND663fQmhaKEkVd5gu/lz8vB
DQuQ/cMz/Cutoelqi+9KSW8eBLSrf50yIfV4PA0D8QQiL0n8OvA+oSdUdotNH82XcW329X2KE2XM
bP1IyE08LM6SSekTr+CQrGEogBJ/cEKX7+aduMQFlLQ78c5kLT0zIOYUSLjxZO4V01yG/k77ms5U
wEJpb9MqnSGjkZvwNiAI7QOogmxvyuh3eBJxXI+1zV5nHQbCTSd4wpokdJbMlx5TUMAHzf9UogAi
hXomozWJNR/5YEOaPZXz3nmQkXMZKUa0A4GxmsvdNwizygYgyImO+z2o8s2Q8GZBldlrbczBzaH1
pxSUTAGZbfPXvGQUGCZYDIRGRJN+0xoeoT3tED7tdOCDb87/mXfT7RfJXoH/ZuHZwaHtXdwSkAHM
syCOVTnyQPBLPvW8R/AbSaV5lL9c4BbaQXAecGchKKH1diPDd33jVnw3vFfOCjLRvQyAW9HOIQ/+
ULciWnYxK0QGZs2uAgMqAAlfHSzWxq4d1Kti0Gj29TR6s2yWfiuEtfSv1MMyw/yBN1IjH+p4ZSmH
ZDKB9vLpb585K96abjhDAn55YC+gJ5WucFGBhEGEJuh1LrCY8ZurR4tEOQ0q1vYDrSc3HtYTLUUs
bOVsjMGvzhOrsXne69fC63QyJdZiQz/jMk/rtd3YT2c3wciyP76hICyRH5Ks1JGQWLxvO4gxoR4F
rxpzrvLt1g8z6gXvi3h8VTshk8qf7n+yTfbdph2MMGWv6WzMC9OYhvRho7+8xpTTOseVzfVy4EA+
ZreaZqyWCsuzdTG0qtHGQ7ZKMdDs8zAiSV2Q0JSHebWhaso6lo/fPy71z7j1uCX3s+YG3OyMgPZH
R39uIQPJLoFFFTBaganr3PZ8iSGcFFqZ182bLzTlKlP128eqoK3SwoAJA8378kWpBaBcSTQ6hJeQ
7joHxAA2Q2nu+JjvQRD6qePvFDwNHvJOFo1jgNgldsksfQL+KIDH/DKRTUyVYzr81FLJDSJpbWXz
0SGySSNc/ROmCoWdR1rQaUpfKThfKLIoYH/yOcPtdXrGOoQ6AMELZ0VUK4tjSFmG4ju99ljKyOdZ
ZIzAspAjq+8ekYeSm0CzCE2eSsG///gygdh56rxkdx6uel/HoFAv8QRKYeaRZPUFMxw9UTGIg370
fg90q1im0Z0EPbjTZ3CrgjxnaMTT2Z6FKCM1T6Vm06DNS24aB/QCjDgtgqY4xzf0W+CxYKqACkSg
P/4w3RKBnijAuhGKlS5iElpm9WxnyWiVWi4b/WYRQ976FzJPBoH4TaR1emPXsesVT2J0nVONocZp
GafPo3bfezoviBO0/MqlveBtv+9JBL9/vJpoE63vdo6t9kIEZIGiWjV44S6tMqYhk191yYeaeBGB
BpYtjINjd4VHeV7SWbwi07j52VG0kKqJsYdPDSCOw6atM+FYWUXfeceufY3HfyQqpEMdOVh3rKBc
W2LOMUwlDI+rUzkGBAh+A3e9AC+WTjlSHlVGqoTgpjVN74CGR9jwsaFc2PKHqeRefe2eOcNcK5LK
Fmyf+Nyjig1TtAMKi42Nre43C5xUidKzGYnvvO/NwjF+Qrp4TJlEgtigolYs1o5CCiCO13Vgugnk
BL9j/Ghy4/BsszMHOnkefX8/JXQyt2+MxSIfMUcihC5Dyx/1L7T3gRb304HwhmRoKPfzOHo0Q8VA
Af+jv8IikqFTleHeuSKPdFDPgPTJc1o7tg8iB2dSK8xzMjMdfgKgX0GpUge/b7nORs13NSM5gEh2
kPLL4tsCM3CV7fn64gJu+GgjOYrdBUltxtL8kiEFM8CNgfV5Tdkp8OV/36uBJjiG5pXNUmhYTh0m
9pUQNC7+Gt2kseiO31CvkTZ1qAwR2DGwn8D9F0o1g1G8MNwLvzuaHb7He9zjZJBlg8EAUwdXzOBH
IH8mtbZ2UosyyEhWyUOqTmikVQ2mgu5cyr3pvq5z3Y0lE0unx6nf65/YPvWsMkr/WrWFegoWcFAb
4OPT8fr2PvChBYqpuO92RbJOO2qGGCUojScW9pXE9vPQaN1dZ56VGdQRAJhrsJhydlQ2wERU6yMM
8g7Y8bX4e2Rr/C7n0gkQKmJ9XYbWjPpEkmF5Ko7s7Xzm/UMnJpgrDU90znKgO8aAA2FBQ4IMFOkh
Y+0JwEUe6CFynHV28jxhIizWej4W3aq1VJj3bkxYi6UM0LtcnOVepfoGxDYcFjsyYFquznfEyDdY
VkzaDRvVPbSclwkOp9iuxfFITRORV9n3MDb7ybQkn3SULRqtHkYu9GJ0gUrZZ4bsnAu1ZiW3R8qa
v0LPd8VRzNUOm/SQC9+4kSTk+8P7SUbP1Z7PKw9P805WPFeut0pOHTTOM2FoaObbvWjHgX9SQhTn
36uxAAlYHXn0nT6p1+/KTDzKJqMnopO7ghAaHE3lpMrwH5eA67NLzIlAvO5iuminxh2rcTDmQI0B
2onM+EwYr4qL6lEnAhhVbw86QBjOVI4udts31RVhITuLUWSn0PDcdCb7OpVDjT31ZL43bnX7DMO+
SNF3i6Qh2BQ+fp2cGCo0J+GL5yvt44Ax5TXdaunc0+kdfuPcQXVnILbFQwKu7sbEg+PmPZYMV4/E
Us+2chtzRcKgVbqJ1sXLtVmENX2cpERS+s53cgYWNLa85OjR/l2Pca1cIfi6BdABuO+DRT3Va1UZ
rzwSeM579R0qFyNVTW3gpbUj5Zacsgw4yX0xOPKUywj7QT2Ty1A1B8ITeOgROzg/KpdnMGd473Tj
uMoxRYVRpx6AadVjZhP2AJ8gcORt+8XS69WgvprS1dSdausJv5RwVWY83CaotYdPmM7+uZf33+e4
mqg+0hfB1VDcG80QNXpQpx9/FQTqLXS6ErD0JEBjlL/TxBRoj70nfM8xVKbpLqIxx1Jax4Uz3WOq
G9xgWEUnisKVF8muKJm4sixLSvJ1MRRpQME4LTtkJ19e/XkxSz9JlHy6gXO038GstVcfayoCKPrd
6F1kWRYr0KbD0CgjMbNjFoIJshumh90oxZ98EhugLYrRZiDo7D1AAMlhXqsc4wfzWGQVFw2ucGu7
QCD+YXPyCPr7vsD/yS9n1Z9bNhJU+9XuULqPAy1UGa77oFvyIbUjbW8YvY4XJmcBTbSxK1lzwgvE
PzhCAesvBk4LtC/1+vnc/WvMPZLIxtWosMgV3FELpnya5K2UFSLdwqB/82in67ughIxXX9NP2WHK
A6X/wIg7KhqbMFfTPiiYtudow6UTU4OXD6HA5Z78B408kxDc9Fh/tF5zZqgiNVoDzq5MfMnu+7Vu
5jRyP3u8rZiktiy2nrUlpE4iDaEetfKVUlyP7ktIJTLcYIyB/KcLkk08pWLKMAz4hGhq8rnMj9aa
hsSb9dCZEPT/z5OjH8xPTEEIRki3SfGBChHR2p6yq6VbSCS6iZcpkCrq1dioAniCqVSDm60FbyRq
mlX3K18Ad/OX5Wpv8x60Cs/lkUtM6QNUn27kpnRvDMiPbPITp8JDk5Y5ZArnOAn7KcKW9bM2SDr4
Q7xyhuU3lSxGWHM2CvfoUnoPjubRettb1RyT/Nvc3CjMMfrPKUTctjqcEyHJca/ToEGdEqhZ2KLY
eMJqg7cY24xd2o6Amzyv2KbItY+kGvb7Zc52GmTJAKkwEjDB9O1hqsE/MaU5ukDzPTl0srNAVfCB
qvvuJXA1LghqYINhie4wh+pU0Tkbx90jdunHkjXvFx8SfMgLb7eJ0L8aYxVEUQyt74IhD1W/gHqL
s3h08YzXLLz7AiNAYzoF/lKSc/K/xGq9nf4d8AxtYms9cDStaoPKQL03RVkBf2N+8FLcsQcALNxa
VDmujXo+ZnyFM2snjsCnVvP0xRbctIx4Ohuw+5u28+IihHYxD/kCWv9lrvdAu8RObqPXBOPyoQbL
Nehp8NUbctC57tlNGysghCfQBlPDUdRy+y1Z8xQgkX/weZjmxL8bOidF/76TrY5Kedbe2SgVc5cr
BZjYYTt/WSKuATMmW8gqim+aA5FwlG7wR5dD4QWuTVVxMSOLTSE0rZUl7ooaJPb4kZk3DmekPd0Q
nJe2bCdrv7Rarb6z0UJ+4kDAh+eg71EegHKfITnQH7Nr+2RLTgF30oVwnqm4t4GfpFPtXBevUzIG
frNTgkiAow37NmNqS4HqoNwEhiJ0L8LiCBvboUQyAmY9fMQ7nRkjqKCTtjmf8VSabSqaq881qwoc
b030SlPjHwEC27nIBitsNares/hHBqYqj8KTw/aw+NAJpQnhsrb8hmBCBHYAugD6Avk4jOdKlw1/
UvlnLxY4Y08CtO5MrI+38SHRtSMjf4HKLRlswL6ZPYruiLg4lHTvjYsEtyR6bEIH1GDkB23HonAN
Nn7nMwwt5L2mKTp1fgT/2EVX03lXUKPCfldu7m6LAWT1OIsWyG8eKyTWYWOSpElhZf3z2I28LaRi
ItXq1hKBEbCsHXopDYs1rosnLku9K5M7vWJHM/Egjv+S2zLNFQBdbC5rvR7CKGjbOjoZnxoPd/yk
/HzwVWDbBQZDj+RnUjAMxWIh/ZTgKK4jnelswfRfrYenlehaAf6Nj1Yas+tlJDVCLKN8wlvrVJAc
GKKwXAq7NFzWABMkgNTFYXnRzWHDAWFynB4ihp2IAqHbswiZGuZLeGI4wpeSWAvJT1dVGfvTmopr
8oJ0uG2M7fmfq0ooI9v5fUqyMuRIPKg9O6Oph+mapfuDwKHXHUp8ak6PBbNUCYKLjJcoq0z2tAup
X7ka8fQ3IdtRaNRTbjirZ5AbJiRiQAQrTECzpdpVa8JZrkIrFRpHllq5a54SClAMp/IuDT+CaUGu
GidHbyD6S/0lrx8W8ljYXX11iKsW0C+6LbTBAOLZ0+fzRmJtuD71hfXnDA9AHcu7INM/Hxq+SiSE
zyn9DLT3FR7H+QvjH3tBqQcwu92bQANhuBFEiXdMOirn2CFIkCnSPZKKwruehncwHHme/g9/Cx74
ICxkgPmsF8qvUVqVRkLBB8Cmn364TobuMXclgXej4xssjBMaqOSUWeX6QJcKZ46VjyIkKirCMvxl
jVQgKyvutT6NY6eOqMcF6+MnxJjf/SYRiB1EKrfDf6SuIGMZkT8TJvXsqE0rtWFQ8PNVIHTzaTd3
uAnU7IN1x3ZAp1pg/rYGS8TnijVpET+pdsuT8mWf6KwiQhUZuVAPG2yPeeQNJ4YHpnJj2Ba8Pai5
UXmUDHsAKu+uAOIOhY9ROfKcfZwawBg4jHcYzA2geEJ9nRQi3bYO3bEZNyCJXbii1NRK23hEkqgT
Yx4B+UCyy5KLHHlBG14y/mlr6FlletDDzOmuPGMcYamkdXOHDAlrCagF0EAs/PHEASZJ3S7D4bVx
7meeAnUbO7DU5Uf639OdjhYv20CgeuJO6i3+SQmR1AByK1NV4CaVZ0UYR3GllCUiyyVBDf4pIdgW
awOyUy5bEsuNUDy2UWzs7hCvwgEBAC2vI393xrBged1+1yhixr+dm8KGReKmj1KDHsHH1FhpsB9R
5pwfRIbNMqdStrrsmwwdmS9Du8vN/EXr/zh1lD/OxjYiL4vG6ZCF8cvIMDgBj2+xUksrTFMrqf26
Lqc5I06v/GBwMTrt0xen+uh+4LKKOMOAflL3uMMawUdhg0SPIGkpnXTev6VZ38BRKj72YMIC3WUP
yIbKYkBbJXu0gQrPFU/J6Y/BEEIsbJVbU4TVLtZ4fjKzmwT9YDyZbQJYlJgNvH711lISW5OaYdwx
eVLHLSMbTVdUnRxlv0FsAX60p5Wrna5wzLZpr9lkV9zY4iH50KbbHlsny9wNZiWvvL+NBFExSGSy
Im05BG5zLFDnLRV9u1FDQb0IJAw1q8F3PVBFiseRhcweFX8CIRCYKeBXL26UpswWo7SwPxzUfNTl
bcI4gNGkW2F77kfJG8S4qV9ekQUYhZPTyaKQyBrUH3eAJvSHenjeeN4Yd7eEFBDX7qfdh+a3OtFL
E5aBx9Cpohwa9w82CMgwdgs65Kw7GyBztrxooqVazl6G3eFSoJtC2iwMbROhXYNJ7dfntcxd4Ojw
WY2lxxAdCy08MC+8+sBF3jIhrCq85YXN8zKNKY67OgDQdG9aXvFgtww4FGcv22sYMvuTvJD65RDL
qR6g7N0qSKNBY62Ia6ncanz8EsF1ACRmdVbIW/44kE/DdEMzTaWlJb5CcYWiRqPpT1npwY7n/NL8
uR8fG5wb/9ezt1vawhQKMSOYsZMvze9v5abuO5vzIDq6ZB0o4Nr+2wEHVJkQ0YVtcqhHGwhyIdp8
9tKHphDo+5LqMtWfoDKu51dHrqfpZ+G7RHRrG3jvOB6HuBS7C4rwgilyuQ0aobgCtRH4m06ljcOS
+/O1MctFEVeQfpuYMa4+ZfQY1lWae/tV9f3GjzHKyh+B/pVqEWkDCWDNVbFLHvNqhCyIJzf1AlJj
7tAGHcZjlMkEsGPA66xW3TbsqF5hRZOMnzrHk1hDHrY0VbW5tXVCLw6zRj+NQc4jMP09o6RDczVw
Jri/KtWfl7i20yY0WPye+3gb7UvEXNDCmdoweQDSRX5zXysmtpZAxUa6h4mkAaT1659uJgcSI6jm
oJUgSLYgZC2VssbyA0kH0vsnORIbmF1Gd6e+10dDmK26OnrGIry8x0WLH5Dgk2va5TIHbuFz0n/u
30AfVqOpaH4fl5nmxlz7J2PuPrUenmm/FO0KKg9NkuverSBBtQXRr93O1VJeglBSsfSyHLwWUgOu
oCTGTx5IFLnn6UKn+cNxjLHC7UZ0eD26umUjM+3LLkSfbV8i2dWL8IOVjYgaBWJU8BJ4QJQRvd2Z
it+BB+MEHaK+RxBo/oXIO26smQfxSpSiZvzKVg4TCh2JAYmDQEmFHN7BAI3vsb0St43gVC/EZckK
EM5b8N8xbtMlEKGnsXuShqGjGhgug2qOErhPSovJij55wR8F98TklpNROBEVTZZrJh78/Pe/lezC
xe1a6boMdhAI66eddkf5SmMp8ekhHMrAXcTDZ7mpnHbRggUmq3kDUh5Na3jQKQWd4izeApXPCyZJ
bJniNPdLxkpevLkXy20Lh82EqzmDH1/31zCabxuGbwg2itB1IHdXsb4i2+ric/MB+5vpH0HdHvct
voX7+cHkOhekXmF+EvCyv3cSgNDgKgTbzuuuSYEdQb/HPr8DxKtnIsMGOG5+D96AHbu+w4y9qejj
mq0pwg9zvkMxh94hZXhOwmCOkFPkMljBrhXEcwOMr/HaEJMGVLoCiRL2RkBcVOVlXhL/1NMNAUVF
O+qWmqGGH3778T9CfLKKmeNd3v9l6Oo77P9Fw2+sMiSzs1Cnc/yVw0ltCfU/oFTyRheP7DS60ufV
GU/KUbUywG1KGNCKXwje1Qnoh/S6K+ga0mGqZ0jaZlcSnIjJCoIblNqgvTfQOntBGFACQdnw+sdt
GxZK46vAm1iRkRb3yNV6cDpSO//+QnAyBTjK87rgMDC9PnQZwVH0JQsEc9SDkaqE+ebr60uf08Ae
pk60VVdEjHRCfG2EaGU2VhOnyK2j0FLpQvkA+WDnS2am8l31QYozrmuujyDcSiSHQh6xG6RXqDzR
1aGqgFsme/R2f++aLoOMC2pTX6C2ODimBkv8U1NuIeWPWwT00WC6WqQmD1e8SgnfhV/SZF0drPaz
pLj0SZqzidz/sj+0I4xuuv6pLXaiDU8UA//W0Mszx2xcf5OCc6MDyBOGK9PN8AWlHRy5XldmnXTM
DZtIKA8W9NYWe7b8MBRXJ5RjyX16DonJtZ59JhtVNJPo1/M8NjVFHiGVa52Dp4O7mSkSovQpyjCa
/6254Ru7bnyBoh0m8NqcsaOyAXwn+q6MIABdjRZzVQbi4GM9vXECtNQLIhYtEAWWHZw7SY9RhRFI
yqG2KsMRlsLOOmDBlYDaz31jYXzYBnYY3xjp/g0vk6+jw/mQGY0go94HBejmCcuKf4u2FQDWfkuz
bYvXw1eYlxCcX9W30SjU/BD5xgt0wYy5gIj9iQGFigzkLGRJ62h/Jh9ZD6tsF7Xz420q/DQgqlSH
8xviY5dUTAV08DmpkGVFgYolz3jew6G1knx11fs/PZthhIdRlmWOwcT0DFkacOoProfww/Xjsvj/
kc30p261bj7q5VG8WBHwnX4SXgSefS+YFNeG9tekNcRDzaQ9Sz34Ej8eDijNSm2gETFMUkhMC0Sf
eBu9yp2enHAhEK6sdAhst4ckI4fEs+KSrquW6/R6WmttT7N6pKYAwZ8b4dy+I9BznCV5ihc6XtqL
KxVSPQCZLMmBcx5qJbvTA2A8cD9YrTv2jaRoWSxCYJFnIV1DXzkgx7FvFb4eBrvOrVHva6QmPnna
zUJT4rgdWWmppCPdGKBtnLPhQVWWk13fJAS6lYfqhns9Ov41Q/vI711jAxqLaZLTKM+S6ucQ5Tmz
as5pMo5IEg6zgD1EzylXu6arntdvsinqGDdXm/mDATtCcNgR/i0+Fa9DLXBQFvVHbNgqZplIseLy
IbBPjV4RPOw3lfprOQNWlSG4QXrUXzkQrzkuYio6SsZwMGb73fX9pxk5Pw41lcszMFq2fVBtii4e
sgs7lPDquqLdZsER05Z0IkQ2q0/jOS7jlBdjMTKuMJbNjmo0nI5lBM/LW5oakXMcNypZUVDILTq6
V0u/+zHoFjzAbp2NKiWCdqTR0wPLvwsfoI+AUXmRisumTgKcoC6i7DNVzrwCjUbzy9Ktv9dZGQzG
5mgVyQFtXkdrY2Sr/ouIjIVSV3F6NY+aBau8Z8dOmbm37Ch3P+Wh1wg3PmW4M0pF9vE16aTPPyCo
0t5pcxhvOxf6UbKb4eGReb4fEEzQcowaRCUcvrFrzuuBCcWAMZrmj/gAl8V1nKGJjeymHn3krLEn
aUCHEOt2dmPT6XsBgF3Od7uI4JAb2L/6Y83RVsA84TCkDf0ffO5tnoqvGmjI7+Ki/gNeVI6JZ7JC
jdV8pM+Kwc3s3KGy+s2IaSkWWgUiOjS1Fw4rRML5HoqX2er0eV43CsPT6/FHYGe+oqN5hCmqxchJ
8a1WWZlw6+fbSTIq1v0X/ovTfzOCCrTKGk9Et8dv7LzXCdaR6W7ZXnbQYfxMKxiGBoNAwVgO/r6v
95RdeCKdS4SbG6Nlm2fnhMJG5iRyMPejzivAwlrF3+tYSXgiF3BcBLcblLpWX9ic0nhuwCHpIo7Y
CjnROMM3v8Jv8hMgI2l6q/naFtatqwDIwsBl3oZ8aNnWWsC3K3fKP0G0/hA7kFydha/FoxUbscoW
BNKozhJpvmRrKbwHkZ1XNVSKtin6fcveQgcdtffU9e5csC7PrU3d6wsP66W8aMei0hpSHkr+LUEn
5+OUFzyYggIw/QFok+MCTOu/rV7DrAgnaeu27xwio8Mrr/3caFE8KWmH5dv8iTKzqfnhFXBqqk5c
9LueZhoXhuhFuySboKvnfMepvIXKbwOtBUAPYJesNMbqxqaQSHe8NZLa8VtM2G5UqPyEEiAwPsvQ
b3opsJ5ac92QYXcfIEJ8Sgo+Dyp1mV+K+hTP+AfliFHmJGznKKuzRt4YEkZR2Kt/I9k/msmwk2x1
/CXV/D5UHsDFeY4dLjdm1zTuQFJeLE8nJAp1xfIP3/DhYXkOygzoDiPwbkbFkDXVJ3jk8r6ZISLr
KzuVf5i6X2o93a44npU8d6uYUxGnV0T0h93PXwQqIcpkM/aGbPbtaImY+dhiAfu6sOF+vRWrNE7q
C+Pb939JRAK62E4tBec8T3+MlW94QSao6fSxKDjSOu6mnBpw4MlHV7946Vjs51CNCbvBOE2w2hG2
JYQcKUwx+w9W/iwC4iW4mR+qjMZXqxqxk5esQs1V5i0ZBfAzFTgNFE77jujz/j20EajnFaUfTuPj
pYDrgS91uaa8KWBlidu2/2+x1GHObQGwE1Sg9h+yoggKmOkbswqK6BO177CWYhbuEbzsFNgPyU2w
SERLjAjbJFjC+qwrx0vmMOwRfaiPBPn6+jU+WxAuRwUmVwOdIc6zlLObg8OMiDZqX6qbR14LS85u
EY5Ljf67v04zo7tsn1alZPz9ees4HB2rPGbPvH/zkFEIWICvRlabLPMHuSD37U0chosN9zrNDIM+
yTeJ7ovynM88gHmvxQDVuwolunJujrowy3Aw457UJobqwFdQdqyGUygOkseaegRfJ5Jrz+OqyXrr
wyIM8XHGo+X9HfYxoaawUJ/bDCD39yQsYiZ4ZMdMXf3JHS0ZJYcAXaPtIifxn8ud07E0kq+QjQWL
xisBIcC9UA1i4nzX0JM0QwsV0rkucVpka4JNOw+4pPu4gF2hv5xta54Qb+4B9TcFXBK1aKmKUP8B
6hzmFjOFiG9e8wB5Kz3TDOMgk7RRDg1MTepAuizp4+urczAG9NK7rY2KQFt/Y3qvHZ4nA8YAKVXt
o+40M2ekMjbqAE6YuT2+aXq4rsFHo+CtUSsUPgXBkVdvLz1yxbI6ZqGKBOhhA2WTlWYV5qfcbWKK
jXH+NRrhcy08hLDV6uGTxsfPai+CA8eTMSdpRXdQ5ddDGHYZpoLBu4lahyqMoqXPhvXcqGfJSj5m
VtYJk1OamPgsliKgDRvKGXTUAEu7WzNAK0hfrCD+LuSVIF1jnWiuqGNwgH9Oumd03oHCVmM5LEDa
uzinjSqL6h86P98LKl1BHH0o2EBYN5wPR31SvglvPuA7JY7GrBM4ZyppLjBcLaLQo4Z3OhO8bGl6
KoHiJpAc4qnLzEMC/NU+Cp/qNis84AQXv/m7987rBurV8SelGqQpshOTJ8YhUZiZJyvyjDOuNeLF
YSdp4Pqhyv7nQ1kLFcKNRKd7B75mWF/53BAiU+Fl1/ePC800VkH98okTe9umye4jvRFJy3rRiZR8
kYrTTq4y+LlICI0yQxRoGa19/a7wYIqopGB42XxiGeO/Rl3YInD2MoOJP3B+zm+MyQdn0j9uL/Nq
K8u5jdZkMlxfr4EiMGQHuUMvceiQKxkE1XrL9OiuRfLLOtt/I0iQMZM/skTM+EMhwqVfCtAZYMsH
HYd8UfMUdZso8bZwKrM5UtnWTifcXncscte70g/6d51KVoIKB0RmwRrrpgkOIxRbHEJydUrZTV50
Kxnf56oVe2m6tbCclmzVydkV8hNfsX0yMt+RZUGxtX/CRBwm+bLyb1jnKJcol9bco/Wbow9M6KA1
iamVK4TdHAkUCF6YoSGLwjh0rIwHQxcaBMuvBUjEZH/vn/rNCwa10hq5eES8gWC9sW2LgYLnLzk5
gN7VOg1KS+vNncgFsash2X9EtUaICzLGiRpQC8K0MqA0aesUyF7yhFpx3GpqYHuNnJiG+qh5CFiW
hJtBrvoNKSrP2ABucYj58qmImtaAdJl/Pgw14wj6xwoXk43QLqGG6oAQBf1koxUuxeUjGpsyHFrE
6iooaBHGLJTsmXYWVG4X265ZB8KvyxDyqIM1IIcSXiVqeXof+7sxOZxRw45zzM8csOelLOOcB8Ss
1Rwta8j5fIJhMRqUdLwhhjbWU/NwV09W6/J3LMBYdLV69pSo5fuoZK0UdCU4HV5tDdKH8fUNsSGx
fUPIDIq5oDtjHCXzdGJWEK5QRmmmMOm2kTA8tJf1uzhRBuVKUg7PA0/2J3skkQGCDcTSuBg7cqle
iczCQ/3WMNpniLn1muoTaY2m8aFA01PoLT10o8iGn2hs94XiwKZPRwyHI3N3xp5/SuUpmtA0Kv62
q+h/IkO0KCOaRsfn1buVrgd67OwSIzP46YLU34Eu+3UYQLTTOETjCq3OP/Q0AV2Aa2CrgpdKyL7B
BFJm8SDNH5DMA6RU7EP6VP6LFRDCk8ghJ3kcQTeh0R37XVDAEp1ofYkFGLPqq3Fmn2BOEo1OFBvP
INVOsfnzvKovggAPH0aSX92vkYJPA4+gp4To3OQwUlXGSQsHAcmkAJ54f07pivtaegyPXODOJ3Jb
/6UPv10Vlmh1jdc9lwIE+E3LHPQCmAXjXIE839G1V+GSdF7kJawxrfogMZKq++F0hcxVNHKbX/UJ
BzNhqoesVj0fl0Ruqsv8uKeEwYHcPovFYYFtj/EwuWtEJOKI3Px/O7G9gum0eoXtNIqxakFozgSM
dRFkC7Vhv4f1aMIGhWhpcJTAk3qS7pGd2sLkGxLE3SrJOwonX8LU1a4qlTEWMR24B0ST+02PDGrS
uJNbO6/IwmWfqwkrN1XJWlJ9bXyGZ5mdj0jaUHfVDodHIEwY3kLnaNnAiBPzh/kJSNv31fuXilGi
mSDasdsVD9+w7VufdstOtAr53oAHVNbvBXpByhUfu9S1grkBEwXGAmV1qTCsfh6/IQ8CowoJ2JER
1ahAXBJ9jZkEkS3K9fhha04hR96nwv7JE3ZVisxgNIGTMRUNszNz4CHf41/cueN42xrK/6+xa28C
rnGjZGSDIu7dabGmKpLgB/HMGq3tNx6rJ9W20BkgLWo40/J/Y3o90taf+fCYf7WV7Mu66+ygX+l4
BWhb2FUrrR26x5qfZ3wnAdfmtDV/siRPLF7G0oyor0aFQy2N6MXhadSBwcbs6f027hl4HAhd1l0A
TS3PTBdBc1ZqylIwrheY8bsHujl8co0ZckAUk2bx0VeB2hzlS4l0dH8CT5Z9qHqTapWKu/gbOUxw
vQp9U6cBLosi6yGkAwpT824PEL5cGb/CczgqLqkE/89W7QFEErbJmqy2SALeieFY67zQDC7izieO
7jI8Tr6wiv6/5kjk00BzXSb2B5+tzoKw4M97oPgzAFD7ozZoqfxMV8hWLycHXn9z4f3AqM5tiD3p
nYUTIuRGNJkFK631RLuAqIsZVjeQCX7rtY68hV3TpX3oq9zIJ0KxxPBAn0C1MFBBDhvXwqv+FAJo
wL4OQ49HbfKOHKTATgSof0Nbj9PNUN7rpXmJyePiC9CstGh43mqC68RUdKMxxmqj7vsxWRR6M0fK
LijSRoJ9L4pO0mRWYM3l9SuP6XLepqKXWG+IP1j4LHnyu/+Omw3qMrZD0kzodsSA/UwQKzuz7krA
wFY3Jl+BasIw7y1KaisGs8WmbLKklR7BW1LfOMlS65xAdrmRDvtaiCI518EFw+uxKrajOSzhfvFL
hINSPlG3Dyp3YA7ta4nBScCWMxf+gp857KhTGqHfdEsyvcOcoPfM0e5kCDc2zKk/K2dJXSyM0Wl9
a15WYMF7D5om9O5XxQVApf8wNbHmBR/SNQXMaUWs9s+Ep7jJC/8iVMXfwzuV+NgRD59Cpuo+Zkss
Kl+yeYUlfHEtQz6jqZifcExC+U3hXlqJJ9VA9Mto4zmA4vmODkNNltmvwN9ljzh7Sp/61be4kpkT
8D3nXhLLxymvstwqPRTXtUXeH0f01wIGOnLxexLIKPcnrggacoOGOmDF9ZQYbB4r2Anm1fXxNVP8
vjzahzQVW97b+rF5Fi3sQCovUYLI67esYeeY4VTad98cK8xppNaoMHe3mbPKrK4QxFKbBYWkP8Aj
cAgoblJuewPYyeVe/qN9+h/XpvS0plvPdqoSTbuNnKMLhqKonfO87OavQ0sBM6m6ip5bxF8/6nc2
V9ljT0+5wE5GwiHq4GKoLSgIcG0WObHBmOS3O7New0RTs7ZtC2r3AU3upNru2I63JSv6EvMYYSt7
Pq2URPjEF6V7jFRqalvxeWdSBVqpIdz1kMUsANEjZrFyp8yiPO8qoIW/MhAIeRl5oIyNTgvdNI+x
k+3Y2RiVd+0qZ2GcrCdwPdvqLPQ3ES0iXknMIgokC0Zo3PEYCL4dYptqJTB9bCTnuYSWRg9xQNSY
OS9E1sojixGaur2ygzcrzrJ2nlrc7RDSojUCBIp3KRQ/DYxuv1YqV8tIx3ePiir4Kg6OObtdofb7
RayuMTiCl0lSclD6ggajZKCGXDiA7huMhX9GEEWYXdsfG+P54FGKIqvVvyGlWKYLCvEKwHGB0slu
plEMg7TX1/8oQaTb7WjdBG7tzMsPH6PnoNeGlgtFgeFcbqVHYAwOiFyovQ/01cDhz08enY0i6OUH
nz3flygF+CFbPztrV+WeALOiOZuMqmvMgeZ2cQT8ypAjPBUYrRtyW5nkmjbb7CVOZCJZjBTEwecv
xuXGmfNwWbt7laeiv8QkjSoWmnVZ0v5vkKpELlkmhAICdDFRV8cbUa77b2whCbkX8b/Ipw+LKjba
ah94kNyPut9vbJv7tOFgpU/KKfkzeOHfPxyJYpVJzoZYdJuOggPPOFiMdsJ7Ig1kphQhN/4RiFcJ
e3F4CnIQ8XnOj2MHw0KXPIEBeUwulbzBcEAzkqmNTdyL9Ams30RhmM4zoW+jHxFO2jo0UyAmpapD
qJI04UqxcEDcHXNFDyYNxY6dSTk1kxfGBhYq3qCLYcJQhvnsEgZ2ACLf01E59Ymf88qPl3rfGLFj
KzXVh0RBnZMUM6DYikw+/qCej6MzcSAG9ljorWTdxDwDc2WXaS6nWTtVuFCJM3QxmSdFMRfSZHhK
m6f0CeYsHv1yetg5BnfoAU5YXf4BR2Gf8v3wo1Ev/ughj4I4N0V4yXLGlsNoLj/9MiQda1IBl95t
DtrRDyuFN1JwfQ9g4NI4qs5KThUfH5oscSRSAa/C5fgI8X7aq34qatXzlhzijB7FNW2aIL114RCl
kch6IdleIGKgNOLytivEIkoYxRLnT+znWrtephQq+PxFY47ktxBoyopH7uyBxjmyDH/Zbbxzikma
xBNFclNlZn8gxVZTEc2kYe77GLOn8QEmUQkF944tay9ALSTbbZkVHm1YKoDiWpwUn5CaCLOhi8oC
oi9H8vlbD3CAoXsfpVaEjndVM2Q/0dtgGTXoS+Qyf6qY2dto06ZS6f0y2w/HXmAGjeBFWdOmWFPr
Evx8Ch7TxTXePjVMQ/TujaWCYtKBtuJuCjGReNSsIjjMS/PdnlOjgQUlYgCjEFA7jbIFpX+tcSED
zowUn1qBz8GNwqOgdA53Eeqgtpw1+lLKCMdkaLWDcP7JjNkXjQU6p7NMNkwzoOEWfeZthbJ0Fr3T
DX35vVY2HzR6gWcsbFmLxR/5TS56OHGnCmQkfYNY9IBQQU8XiTWWGdyGtQqvx73+aGw8Smpv/P/O
qsxo4fznsZbMErGiVWij0wYy2rcJ0kH/2mB9Oadyt6VKIxFLP09p0NM521alOHZBIeB/iGONxBqr
AVlec5E7Tootrkz7fEiO3g5YTA11DmNXu4zeo+FqvITIbZ4EUbwaaoAa2K5dDyh78Ubpaj745N1S
WZ3IWxZhK8c+2aE4NnBWP8LMVz0nB0mageFl2VF1dqESLtI1JBRX3XxPytiqH0cgZwer3zyCC10p
C5UEC+mqYjRbdWgcQjgCZQr8cgxNYjOB22kZJiP0uYDNdZCcFHTjRjCDbtrsckjVEHjFGUxFCdGM
N9JXkDl2P+2jDFYGreuVR1mYLTCT1w1viqbFMQ4bOGg9GmvbFfaaqVZfgGtA7FIumqX7xLfj4MlK
Txz1F7+WUr/+5pSWs2ZUy/HHbnzwKnjZ7XgqJJARh6rR9usTZ3fpZ+UVrv1eM6SCMu4/hIr9qjlt
Iwbi08WjlgIFz6uB+UMc95rvLWZn/1b5gx0VzerSEo8isvIyO85FSe2ZyBpuOQAoyZG4e2AQKXXa
UIv4MBT0aFNIx0SqPkLPvLMcudulwVhMxNaf6tlghFhzy9Mr8sbKEc16L4PHCMobPLrRk+eRCxYM
x4G7/JMrjVKUog5Qss42hBeLwN+oNI4kmkaDemHYIsmDjldwWcxIAzMRsUOD/SeWRPGQUF1iCfmB
7Kdo/RL4jyQtOnpsLOr8V9YtO/886RltPnkY0IEeyR/WaoQiT0/54hDDSu8sjAA4w839UaIER026
OxOqyQzyrXdOEQV46cTtMOfh9l/de6IgaDGjI4ry0sUOH8IVvnKzqfXUvhM5HnKdQotsDr8WZCYJ
HwVSjgC2RwsQ1COKhH+ojC/G6gLSJhSFnV8TLr0L4yYe+9YIXYN6eTDjH8jP88twAStKAn+WMnBp
R4ieLYyYDNpv/QVsN3XXa61BaTgn0cz1fdqm11+zetFOyhYSi2qpKa46y0GhjmZPQYpKIrXwsdZv
YlMaw07xNQg1t1BagE6bmZOHdAWuvf9Rl3Zf8BVcihna0UkT1BSuSFqIPchbKOK3cfiNsst4P3y9
EjxWW4dfEw8Fayug3DavHkMQQQj3uUDsPGVyJQvom2RASHKpIWjwzmHn6gLaqau520QH9Ue+07Rc
pCj1NiMc4JQFW36TvU8cx6xvrrgDpIoeDvsVVtmz1qc/r2iyP9Sa9XM0nG6VqbljJ0W4b/VhPO9W
bO9dU87w54JZHQTEILMHb3rPxmJWoK6VE/ldi8Ryz5xtFEc+/jSTtal1Zb8Wo76TE7MhwC86pMvb
lMPBzk8b6wtmi/8DflAe5BHJTgQjsm3nQse5UytvaM/LXdwj9qowT+9qHhAp5z1iNiMnSYMVVKSN
HNpp6u4tG1i3ebylfhhGspWDPIeexPPFdko/l3bNQhUXCSVQmi4c3Bw0LSzuBqypiIJuWdwBio30
RoPeNzPoW6ezp3oWeoRx+8nMVFt7gnxpqWeKpK1E0QV3fCASFPv8q+E8A5y5U3Kah5fE/3yOjAEG
gXC2YVJXUDQStDLJT56NIl1dyXnAtmuGFhuxcYsTPNzbP9QaStkkvl2QXck/YG1fJN87+r+j/zyp
DptEvhbfZ+h8vEV21AyzH+d6n/VCc75GJhCriYNApTsNBMfg+/A4OqlZ8j+Z5dHe4giF1LWkANi3
IEX36uMT1kPeXwqU/9uML7iTBQZIxMi5agFSE/I3x2jAylwj+hYY02dcDQmePfvD0yDIGjbwE9p5
Y7VAso6KSSVIC5+Rl4ZyyZ7b/HI1Df3rwH3E5cQALFnBjBYqVAtuAJrBprq1bX1VvyltLRypmAOq
5g4/QrYlXQFaFYSCr5dYxNoptu14EMtWJA2uteR9jXPD7ATrINbNNgm43vmApMh1neexlU73aGue
JTpYupuArFra1/C2H/5kxn1JFmfSG8jhSR5gc1OcF8HKat+IdN1zj5H0sgURr5XDqfSl1N5RkrkQ
Yh827S8va8vbKrSWVmUxVgEQ5KAZ0P7+exkXayZ5iiRGUsRf83j+oV556hhy3Bkd379/EKl87vT9
w57upjd2Ebol/Y/KfgFMW9uS8GyWaLVukxgprmXLuh9ZeHdcwG7BNxPXXCLzq3jBkmuglO4geUWd
wKTMA+pFvBrB+m9IGcDVrWYiIE1tvtxMw8OHw/+1rve1Ex/uv0+IyrVTrl0sC7kQTMZAFhq6Ptqv
Olmx3wQaxkvU9uhSCxVtmmPYLJKyK3Eb8h+G91BNqVGZu9CsziI5vYB4bxVM1Puj11YMXQnoxSNL
nMC1+g4SbReaskdLe0y6egxldJTGxeajKHrEr2pOCnHKGZNGlz1RCJzoxp0iT6NnrFGY/Lv23U07
H3tXA/wZ8Ci1vZAvAogzUcbg1RRxIGIHZv7KWke4tCOovgjUs3X0hhYIVvhU2fu0EygFVrLoyAXl
HtlWjJ3lxjImroBfhN/I6rN4eG+07RoxOhWos3SXJFhltRLGTfWNgPclI1IusBBF7PseHTVCud2Y
guQNM18xnrP8LnhqKkyxCSJKCV0Dw7Yv0wvirBxa9ehSvHc07ahJwj2ArsVB6mkmO/5XG3LKk25U
3bA8wyGZlQBjwbUp1k/v5KWkQ7UC8ltvz9CVe+taoiFw0UZ0sNjh1Qfu3vRvnt11hijVTzlq7i0e
jDAU9OD4Dt4lk74kpKglSy4YY3ncfQdlWzFMTc69Fq/UA5Ow6BTZcvu8/umaeV/s1g0NiSDI7iqS
AfzOtz5+RmONydduwzhjl0scDliPVM4OIqqllICPJBgILRET0EZOwTChTWzITUhr1DfKrJyJnUhC
yJrxQaHGrc/FJlKpIbdSNKyiFFWHLXVJpPKgr3lWZ1/gjiMkO00Rh6HclSWfee5iakSO0XG0MsAT
aIabGTUNp4G18fL09B+QCDNkdO1ia8n3nY7kn4dDiN6mqFkcUTkUJgC4JsVcCDpIZkbYeTo4RFt5
JWJUCvPQrcgG5KZ0HC78I58xIj503lVTLGExLNYA/qsfrJoXgW9VjoQj0nl/MjVBhuFsgbG5Ym4O
4ky4gL0NbW883wqO5k03wtiMKX+kVmUUbQRXsS9DR6I2uMpew7Y8dLM+bsony3E1mtAzhM4MSSrx
CpkQKfib2H3gYBtZpYVCH6fpfLveg56WX39GgUUzOsYQ8FgyaG22vY8+bPFQWKFHKgLaF3cluK99
NXkKes2eblazliRJaZCXCCvvD2Y+MlZjQ2RIdmhj15enPmr1XIgYDbSaqOJWSdoHt3in8jtc0tQ2
sHLQ7I9pm7OoehmbxnA40xRgkLGUbKbT3hmH5yD1XUBl1OS0K+WbL1RmfA8JdD/z+od7/42reuJF
UyxBzcvZPSkK/CNz1x9MiyoN8m2H8W/Fb/YYSPw2VYVX9iLpo7+7wUNW75LAjYPTbr70SV8pliqa
Jp7CldWLQP5Dm+Saxy55DYW9oCJek6dwcNv1Ukq7K61bgwChHFfG9sujqbXpSSWpPuUwkUW+HYED
QVnNsRcRxwhvSvjKM5fMo+L/FJcGCU5Eo+9Fv5DSPEOu7/500iVS2AOlrahG2bMXiT0f9Rhd46L8
p9R+8Kyxl9xqYzJEuk5MLA6wVbo2oLs96pka909JxvuGg47+lytRPm8iw4mUFJsA9Lk6QiS3EbHV
3Q+MaJpdOV5jWVNv9524xc56vsUAI2yQ1PPx3GiVFmnSvBzcaH45WFNKhX3efQC6/TpxIRJ/3XUi
QLxknfiL3ju6SzFqEV13/n5YVOJsJCcVMH41dNAuFst1ldhPMHQz5sNtOYFsyPsITyxfpznK4wT5
ge87k+ghfpc63wI16R3jAEhFfS9MudixK6hw/VuTTzn3ukuCSNTjyOw3st6nf+JtylCHc+pQ0kGz
TqPzpwQ6W6S5vI8vm5HUTGUF6X28CNu5ZD41wuC+Ygac1yQrLG8HOERfm/joaVTEPovDP8HLysyi
QRyWbjz2ntZ8vB1NLlTWVJCkCq02cSONl9VDhJ3g5BvAtkPHjMmfbfHUJW9z/gUkyWd+b8PAa2Ob
zyTQHxbszBL2h9SiYUcWmI/rLeFGnEJiiq3ymTl1PtPMPoAZg1nk66eTdazlQCo1jferzYuFexcF
rfD1d4hMbAM+zOSNchSMSbYcCsH2uIEfsGXv7sHs5IEV4xkfSPXYmxKxvBpCk177oRVcEHNCdFbU
qVXOKGyzOFRY2Fkc7T6d+nK075vEZKa/U+4SNLckcZG/6fBSxoMqKrmaP2uCc6aQ1FtNBq/1qdc0
1zKuDeONE5kOzRmtEx0gM5ZJ25kvWW44mozNYiVjmi3pxOZEkHWi7EZLmCJ0D1Io7og75qxiEniO
orNba+8i5Wj6zmus0+/lcziIGP+lqEllChvqoc1xidmejtPaoltlAP4U0tJRvvNvlmq20cWmeJ8I
5+Zw/ANmmXFCBuP7nGLFfGvTL6hhjOxrOr3rQlQZ3ld8/WvOs4UxqYB1FmuTdrN2fByX696ra3YW
uJzz+jtyNdOf7s0NT7mBR3/wTunjnqLcm6ui2yswld+J/BgL/jqSl3hw8cGe193vILCVU7u2Eg2N
V0vrtpAWoBie7JXJtURFWQHp4iRiyETMJnK5A4fdewpKCxrTXVnMyiCaAWAMjI1oydVlB6dGw+Q2
9UtBRtEm4ThHIYTr8jUVX7cjbvxg98mh47wABNtdo79YaI21FBQIgETKHnSSWLyq+HcKAQ5Mv8/q
t1Vk1YMCLN5TvYzmL2/dCAh++cPhNaXgCSkJMzoHE750Kv/BLz7cnsxWaEyhjxDX4CmeNbNKBqVh
3o19GPyaoD9puEASyPOvvC81eK863N6RNMgGp2MZgrvbuzockEgRyEpjzEWIMSEzH+f4q/Urtk2i
680olOeWU/w1hl4Bh+y6cZfKighCOUu0NRFIc3Pr8aApwRNIF2vIFHJCJTUQJj2ODW4HJzGEcEbF
yhYhIktqyg9l/o3WeDLfKZslQMWIoo0QvqZVR+zFnr2zgRqW19QXLcudjP9/xjarUMsum3TMhRt5
9mH5JR9YnOr74zBaYaJaqto4yVZnFeCKlbs5Ip3LhgyP8oCSUqPFqPyFOhTSPcsNQHIxBiRfW9KS
BdjFu8cb3ZhubCCi/wdH49ia6MXXA8wKTKCa+YVTPIqQcQ7w5InpVPpZI2xccEX6ybUDwfmdrGoc
enyvOxwwI/Yleslp8ygK01g3MWUysrntyfcPKSTJJDyE/mVxCQ3JkvZbfEiK0HUAhK0ysPqxoENa
2HbwqYQSkf/wuFwxWAtpOFW2W+ilqHmzvaMLQ4BMhWJ0AEIHOes/71SjHYFHqkzwKmZpFKJlijlI
x1xJiR6G6MDNR5e6UundqUfghYVU70REgIehbW9YMrYPazQcJ+7H0yI1xn33Qcbo/odYTPtrJbc3
L7tWXRbudBEQKptVzeZ8F7lFHnpwr+VnBhK7ZYeWbnbLRcQosn+y69/oHp2+Zlindza3HfZllzKb
18HF0s6L84U6r6xfrFj+Ear1rBsD4rh18m++5Oe7Qj1FVE6IkRPF81M6wnINhmmXcZpeU7ENK4uX
RrFIqdsbKvRm+0AvY+YAQRwmHlU9WJY/tVPgWVJMa7iFwn+St4Q89c1V6hnHd8T2AVKDAlRZ7h25
xP2qDeuqtfIU3YLPfW07b4OEt3+Nzl9PLA94KWJH7e8fVx2XUtlrzXVs7GW52mN6o5ng2sHBs12w
3lHQyLriZmFiQ4eNLQ4uuCLo+AFUjwafNC5ypGUlHO+DMQQoK7ZX2lXu8jtBmRaocR8TfqpkVHVt
2NhOrVCs+KR1DaAgn5g7ejtZ23nsBr2vAdEJVbmDY2x1GAlvKNpAvC51VyUGiO5f9WK8f5SwFiDb
jtNee48x5AroerL95ci3r3HLA2dRYd20XoZzR1rdmOFBuXcz+l7jTNofNl4bYw/JwWXI7VBxcy4t
mK9v0iZ+IiyJwMXQIA8C7DPb7txJ5g1a4fXa830DvyZPnlniWaR1CAiD6l/S123Ktc+szM1d2ERb
1VN3M5zvns21SO6xzVRmdR6xmq7HyBEte3/SeuoNHe0Q9Esrb7aQGXCLtJHZ7+BeDUCx9OYQ4W4g
+IuMPjsNDSqRgGi5loVBxcNrQynq9xHC82pMzbmJkr+AwYqVd+f0I9iEDgEprlJSkKeuo3QxPMZ1
stl6WLg4XJhNN08cCIIRTdQVMfRSn/UhC9US7PWFlgNz0hHGleKmhJMLt9iBty9I9MeZ8U5B4+jQ
Mnvp0y+uLnUK7sh1gZZhI9kijSTRqANPHuJOe43qT9i12hd3Kv88IpQvQrjMRA20KeKX5xK78rGZ
SCKcxq1YrEoINq/ZW0dLkIWWbmE0yNf9GZtQPhh5ZVWxr8fiX2OOtWJH9q1yt8z2e+vUzSK7D92K
hKzl4gELFgN9BPGjOXgpK0S1r4Yy88BGfGkcID7+OTTm6xanYAmqRDTmDjkdXCgHvAAXT5ZtzCA1
xXMtQWPrqRph99agtyv6Q/Ke9s2bvw+Ym2baeMTzMa57p+gPZPqomzff+0VbEO6t6VeG6SXVGUS8
4BmtMdmQSwlsCgRMwIe6T20K5nZhG2sLTc5GL+7vF7dCjhIRB6q5eHrhyx/e42MJO8hofQHB/kc/
9/s7rfqCcp3pHcBvRhqUcmYv18Nk4GZs/voLAXcuHxwIivBrDVxjubbZixhCGhxwrHmGsVYRz34b
opsyG9/z/4icRBrjV7Dz8xs0g0xOjatg2TcfH3YkPRnXBLSWGK5DYYldIEtJRTLb42DPCD/6XvfU
iRV/ePUjw82Y/+SLqIu+AhkhBiWGyor9EZlBrIV5K6kU3dIgzXCTLRNrohfZ57mJq2oEc5vOmuqf
q9C4nauJNfUOtH+CT45kfsHKlY0bURegrRZDaJ7BXC6r0sE1sPSDFrVdsSS/6Xf0Ff7Zs2Oted+U
at90rSOpIu5x2rVKGguoulR1Q9Ydyjsg2KQ/DnrMKSRXFnWQ+DYvp0yAtZtrAGxOnx3Fxrnq17SA
UwHj0vPJppPJvsYe+RosrtV9wQl0oX+kMlY+lnbxAP/5ROeh0iC3DKc3b83btyPFnBixh+G+xzWJ
qFhlXzz6t5hB38S6ZsLcTRZPVyUBngj5zcUOj9Pdik4ZA0cNzshomywX19WwzFoTU5T7nR9jMD/M
T9KJxVKGky63anN692telrjBrREAGs5Xgt0H6oSCYuuJhCzg6UkE0BDF3pJh70wK7ltQVCp8a9Dw
bU0EzwuVJgHaQVES1Ym2pDxE6P6CaErjr11AMpgKpYaehqWq47cqBKvtxSHuFx35SsjW9xkks91y
/cUE6Z973D4DX06THFAb76/sKchZMO+1e0/xIbLvCarX16hXxqcwdOBSrn2tXJ4GxrevXrn908BM
PCoPz3ihhI66IWAo31P00OTW6e0S3mvP4gRGhkqAaZfAOF4eVY6zNyyyKcOqb0Pb3G1Y3DKGeSvd
/Ai555BFfNf4A43tIgoMac8F85/6MbjL0Qmmyg2PZWzDa9y0zrDqwpCt+qds5m92AEGARi+OuZVS
X+xiY6W+stRF2zaw39DByGo/F2MSW0hDF4l3sMFDPqrkxLqUAFe2NGIJe8EacEtCss7u3hgz80Gf
vHzr0jHvjvQEcf5Zx8ZefOi4UzjZlGMT8DZHEU1tiAY3F2Dh2DOSqXjEPx0FJ55KfFYkpSf9kGqX
X2HOpzoiZHkBmw5Q4TcrH235iOcUbXk3OmJfjqDLW0oVpuKxUGjhxHigKU0DVrSxxjKtEpon2Ohd
wFj5Nu+gevPWAtOcfqbKYR7EzQYX5iZuVgzyKBkqltu4AJIWh/ao43P6oVQjL2ImOpjXvGMLCkdn
To7OBhkj2WlGQgbq0tEXCyjk2dtiSqS3tGdw6Z2+VtWj+TRg3I8ov8hoRM0sPqE3OSiyl/GSMADV
PdsKHOb4XbPP+Fj5FT76wv4L4lzaLUm2Y8v/GpHNGwXP8nvM90CYCxzIHHaIC759+TFcpodQMrkw
2hxIQzTJ0c6GxmiMTldhmhAmVFCiYr4q8ujCNn2GYJAgmPlJe0mCoLkC5Qi41VftELHwKhQurNCL
fZEfUrVNaVMfpAlqQmxIOhTVk5J7wQgSFkFmf3bVhaJDeKbcN4vtWJ8AuVFDjWk1as2bSf9EzOA3
D+zkiWE9kkKldx8pNdPFx5aIWdARS6/o7XeNosvMZ0E8gckC+BrVtyc7B1U9eNff8eK4gjuEzNTr
l3V6N2ctyW+KBA6jht5lisCxc6yR7N3j56fI1t1whgfJQniUVpH7ztwoyL43BXBw1JFMEAhvg9bS
j0Mg2QCKn2ccLcbH9ZKOuLB+a2hHzxTczXJY2+D3Dpna0WEc4bARgBWhLO18wdEoAI4y9auNDwOX
TK+j16MTiunV9yfwOfHLfk0oh3Xv75roB3ZGD3D+Eb9T9zyDZE8Dw8Ua7eJkFPcxgn83wa4EY5dn
Zymzwuy7LxG0t0Ae9236xqZjd97yO6G/rpHprdFUUOn4wQs42MhsXNOOOA1cVXJ2nZHQIqasBS8u
LjFpXe26nM+nmjFjK5Rhmtbnj9DCUv7r1Z1FSELQXtgc3JoxO6TLEca/oerYZ8MWlovDf3yZ78Q+
jcxunqiINm87oK8On5tTAlBMMfykH0UcC7Gaaio6SiBl/yD6byZgfF1Ak4/amJR22R2YBbdYJZqm
+Irtnnqz1KS0et1cHUwZV8YEQlCT4Y9fl8WB1e6do4alwShYqbIOH+B1/XvlYB2zIY6LMPqKXlZ1
xUjy3I5gkiemc/MbOBxPzv9XShGfflhzaDxqXCak0vo7yIrGoUJuyDMjdJ+92NGebAKhobpxZNvB
N261Oq3IdozoBd2rVkIF5fX8xrCtEhAzVTXQMueRjAO7HyQrovWIgu/C5ojj56/RuXgyFTQSE+IC
Qb2AJfnlQJEAIJXs1ccoDT09igxjqICWk2EwfmcqZHpZMjcLTc6y3/a2P95g5mb328jnIHwnbVV3
nCnxgZzXyMihwAtKG9dGl65F4ba8YT38g//kbRxO39zHCp0gj8VnQHO+xj8CSQHPFNMeBAHw52ex
fwoZ660c2M/Te1TjryQeshGoczFIGUMzi1ppEGcYT3yVZJp9cAck80l4B+i2300x1cYT53uP7039
cAVNOMR3Q/+1xkGVXmUOmV6JvwzgUJtpxRD3HW3n0Uuw1MlirI+RCH9PG5fpgOTTq3h7Xw6UhiGf
dnrsuTVyIm8WZQVCZxe9T3qVzEB7pnbypGyOLjjreKygtqf07+HtBMLMaCy41sCfyrc0wkbq812c
1crzWFg9R2vJ+84qz2w0S3/SltztsviO/v4rY5IL+2F5ZezVC4OCoKtsW53E3AFi4oTOJ3ywDHe/
c7+B7H8b/mcPPGVstpZOZyHe6eFSUMcJr0QwPEZJlop3g/4iFYLzgWthv9LvHAoYdi5EBFAHoQH0
lRRJHFrXFlVTfXOm4l6iP2ef7Nkeq61SGqNINGtOPx0G1m2m/+h9kjTIxaWvsB+IW6GCLkTPwXcP
EfS1hDmGxf7v39vRhgc15Am5HX0WS8ps6DwmaKMfSRQIeiPx7ohGWbLlKceK2bnmAx4eDgwmcBy9
sM1NCmj7mxa7ZJipcStwkzUIz4L2xHpmztpEWOUWBjNbfgeAmmd9B7bFR4du+tFHHozGuq5bSWPo
gzmcinsCmQSsiXiza3/TSnNUoXeufsC5f/Fr8gm9fGopYlRuTGjSjJY9D3NCVIuNQyODq73Re1UG
53SdRidTEW1zaKXaJrfz6CzQit40FY5HcKN+32hQ86aOpRrV7TJQaA6Qp4NVyT6JQEMQDkvKeZEW
cDtzL6NkC389C5XeMuokgx3SPLeHkF2N56OL4HNx1Hx/fk9O4Yg7AgdbdU7ooBLfdLj4eevuQ5H4
3y3yXnaJJKoYziMI7ALtEat8FCOLKM4gHcDY4Y+Kq/LFQUNcEBDk4mYfIkdK9h+yzrWO4mLt2IPq
J7akg30+iaLG2Wc2925NxHa6Hj6zccbfZchWr/bMairXHlDfdM0LYASIzPU1dOcWrB+X+WhZZLKS
gofP6dcPgiFLHra2iU71S6Euss1VHf0St+T0T3TqQRlVF9rWCzD++V8KE7DpOpEw+tcEZDO0B5l1
sYymKILrYZBV9XQI/BDPCF0sa9f98pnZEkTvu9stcaqciupk51rtXdFOt4hlZiMcVGsVYWq04JGD
TvUVROVr+wRvONnd5wp1l0osgrMdsVamMx/IZDN/XKuHP4jBdu63DVoiEcmhIvVaKExC1JOFq1qg
zmJ1X0BC6Ebk2Vtan095uh6W0rSvMDyIHF/a/6WQ+qSPCid4LkrqWk5Rr7gtvoKiirASyc6CA+xw
1fNP0GDbOq0nyzPfJ8HJW7H3b3kzwt59kND/uJVOItCSQzP9ZNhfbEaduoKuEa8jLsqDfqtdFrNJ
wtxrQMbCBctMHGmZQPtJJUKI9UwIPc8GEV513WUV48uOubKIoROLIECCc2BWvw2obI3g6gGgxKrz
82HV9ZJKTUXMPx+q7CQ97U0qZdm1EEYmlsgGGoKW9ptYqLNeq3eiuomOQDr4Q3YYFUg/kwYK/cVJ
3KDPLGletUwgaL70H7urPuyRFz3fCYu6+X0b14SVyA1cVCetOH0Fx10IPgVigtQLoxvvv0ikcGMd
FjQ/i3QnYp+CnmiA6qFl7W6ZH3C6lbqIbsX3w9vq9pOmhk6CIlZiZDMa5f6Fx/+3NcE/LgkSHEnG
kwlokHazFM9okqNi0IoyLgS+EatV3SRdnkI+z09sy1MPHOUDXIC3WxT2A500H+eAdiEwEceWP2af
wmML567DM3VxKKCu5LHNbDn3Fault/Ct7hylHKjj9OB/SBE3/Yl1qAX11KZ2y682UmMevTubLR5N
EzvPfOHiqfkowKpdGW4+OlVmH2tC1hJ2DYzJi/he2LSxjYbrFUtSoS8iBd3sQ93QjxHCyakrAhf8
1nuiTI9n2ZST/TgYZX1Y3VsG5SrrIGEqeEqObs7pDeHBSvU1wDI4vaiNkft6Xe94BbyOdZryFM6U
34tbYW1qRfsQzt1/q3Imm8csBKtr0GJ/YJKmypJrIgTGCpPC+fTyux3215puhjEbwO/EvCJsJ7zr
C2i/pPEfAdiRVDzHnkrcXN3zE1ToINBPHD2x/x7/P49NKI7QD4OEQM8XrurCXQaz++DgkkLm/gar
k44Nrd5R8uNn94FyVVijSe8Zg7V5SSpMkoH0bPGVk6eMVQ+myFNCJbPhlq6tAhfwJGbXfwO2nAtx
C4j6K170UOOVY05M3hgrv1bo+1464BqmX1JCFtbEfR1NBM5R5JSm5Ez7FO/w8JPJUoL849MCcXNr
kqmXGcR4ZcbJIHT1FrPwKg09p9IeuI2hejjPK8ZEG/P4X2X7dWPweY4kxbf5QRJfRxfv3aj879hC
C9U8zMgL4EdurRtJO0em0yttDJ0oznEJ9/fZ/w2SN5PH/7bzFQn/rbzlw1pLC4YvW2dEz6UK2Hb+
nWwbM8I7ROCz0XAtm5kRbg/eybY1bvFHPzulNP3Rjxc19w32Nz//HQdT/2f2iUfFUL+Im34qeVJ/
tI27xux6SXYtgVwbe0wAioFCwa7GBRpdycvlgsSFrHcyfhOo2kGkchNosFgWD6p+nHRUBeTiW7xY
eYt/49efhvaUEKrV8Cgmg0a8+zjyQBz9nq0rMc+IA8kyr4m8He7bwKaN7d2l7xdr+ULOgPRRsqF0
OasWM4PHNET9PsplpXWTQu8nFcK/liqs0T4yXtfyfyHFgX8JrZR53H4vEZ3EJcViXZEddyewv3we
YqzHC11OTrAJmuDp5zkaNzgDDodY5W7GSMjS51dzPPvvA2KhCX8s+fOGT05lUZRrq1kZVFADa7kJ
VFW5xeZdMqDaxYyRr5FgGui8h4G0jCbnAfnaRrPndDW/ESce54fJ4vev8H7w+xCxnBaRfXtMIKS4
i8f9olxONGDCFKkGH7Feo+VVVRkBMnBqwTsK5WHL9YZy5BRNf9GF9YYAkWo+JPj46mZTJYH/I4nD
XadU6X7lTBtewpaFO09aYOY2mmkmDVyy0YwQzW5mJpfdHt69Key5Bz5AIMXuZhItgQdcN/IPIDnS
Rnug31uuOXBgD761lr52YXkcztWEnwfpYqc9QGo4HqDS2QmGcSrfaHH6sSyUlSsfZt91J45rmXKP
785F1NbaD6M+j4Sys4JdMBjL0S2EVPmHJUAn/TXUtcxglzWAfSgfJNmnDMrQoGHClNt111WY9pKT
3dCI9LBzgqPp6bMrUehR+dKzp8TxGjkwPpyx/b62OWVLbykNqKZHHVvKGIXpXFANqjAweO1rSnS8
KRB+oiKf4lGe/GOPqth/rY1mOOqSgxX0HtizBthYl1gtJVvJ3yuR/IDBeWlre1EUI2BAZfE5H/HM
auTyTmJgvG0vE6VUN/zg1kkNuVbdaLl5Ig3MvK2uzJjcnXxGiVLlf4y/W/QT26fac25o5Fn2J72W
qU5JJ5mbzfa2LkZ/GVAjwqwe+h9qG50dcB/GOr2p2KWTUCS2b8AC/Yj4tskjr5sN9Kh7202eTflt
GvDPrE5ywIYNMTLpMZz3VQKqLMMo9yCm4ooWMZJLw1MHDnTdezAratgmFEOs7iDbA5fhW4weLleW
+z9+mniIBCM4Jz77SJrlZ74jd15974Pct32yhu+DYaOCe7gxH6iDd8OqAPA8yNRK9UKUPc13ZF3O
Nqt4KrMz0xMFMdIenDA5ZuhioXZKp9TG50ZyaG053YmeozwuaIpdRxupliYXG/VSPyrqmFOgsFYw
zh5blcR0eg12bX0OlwgcOtQYJfUranrjEgoT3N91/Ap2vSb+p0hRgJuUISRrPngOO7awG8muacYI
iehJyP/iX0/nV6wHtCfa9PCiQIbbb71LOCTxm4p2F6AekR9/meNO/ox4N78ddKSfAzYAh0r9DyRs
VkuCaYjVpM9VIWrATuVJFCtBu6F/N+9b0YAmUsDqeex8GgcOy6QKDnA4LK8TUfkh3EJ+nNO8Ckka
IZcpvYOCnv2MNzrxG4DW5M5Cu5qoI/jYBtjWzgbSjNDHcYzXej+zKCIVrGVRYEL5TEIqprb46hhZ
5T2oY5Qb68VkDH7cUmYX41cxO3g+nUzzwItZmgXh8mw6a7IzmnqsMT8Q2bNjChYQj0+jmOKkqrY4
IGqhAZUxsiu1GlZlYKdQR1vxolXnH4tTQeqPeoPz2RBTs0DwTRzLMC+SKZLZaThC2uoF2iSLJbcA
woXKKisRPfVQBGzDwuwTQyo07UmGpUo/DINEO5jL86gORu/wWW93eBIkGnvj1hrnzvn1KVVAYvDH
2SF7WNkJqy2vVK9KQn+kVDFzTUOWMu7c9FtNphMMQSyb9xa+HPV+1ykgUhhQ1m8yXXrAana0dzqZ
EWvLQTx1NxuPN43weAdgqkbnTH9pn6WmdaYwWp4HHdRiknO+K7DlrUMNf+oVbPDBCNFYQmJl7U2M
AkggNLRJnNOMMfMWXE/ielkwC9mnv+ujhXd+qHfOD9CPvdoyhcdG5zR8A9u1IgVeE1acGC7hRgEu
vWChSBZtcB0FuV98HN/uyE686lOqGpVKaKlPoPdAV8/PQmNa84kPKFi/uJlcRHZxAU4agaEXOob7
/omzJkVJBPB5Y820GGo4SWb7czGiP/7Cquw0Qp+MEngNuyPLfruArye7OzDRxlm1jINWusjmJrUa
0DeMM6fCy5o2ZIPALKAK9JhSBa1BVCSDDNTEYMdKLvv9El+JnA0XwpSV9wP6sXeosAk38bTtkrNw
Q+7WyPQdw3XqH8TI3cPepvTs050ywxXGr+ikz2oWB6Ncj+20jWMR3npH4LosWPPLsA9iVaIKscFl
YFW5PgpHNiNTl5l/ByZL7Xa65Wykw+h9mjxb1d4z+8RmjWegmP8wFxk7q0wqkRVJ5iarZw4KePsb
tSlfmzaEpiDMVoro/jIbwgMjVQ3g749DMj0dc9wy0AWW2cKMK1uwnWm844wIc47ySz0abauZ4ow2
oAoht7CuypBmQZYN8y3AjQ/XNLU+9w2o+D9p6HIRpMaTfGPC890jBIHucw1ksIjfNUYFmqSySLcG
tMzQBBxbhrUxQ15cgO1FYCZI2bGI+EELeZ1zUTLxibRbPM7vImEkreyn+pf+kp18++LF8Rz8ok8J
lxbWmVA1gr9nJZV0cK7YD2atGcn5O+swlSDTzzjyi0p5QM2SY6J85cwC+Wh1qqV4ya9ivmW460cg
npvDBfsyqB69z2FEAiq3iJmlmv3UeAyluLOyLcb5go+bwNSi4VBEwBBBadp+gc+Qow+txcBVHDs2
qh9LRB7LqUwGWXexkDcIymH2msXmHZkD7IlaALF8Ogl27XV2kpLnnBmWNfstODS2MJ83BTdKl2wJ
MQlYh167VxRV6/0AgxNGki4lXRvG2ga5zs6B8j6hERngQWdeYBFdGYAI7VWNNFZBcwKVKSnvqAF3
oOwJbnB6+9RPk7DA9MOv1TY8Ufhep4+8vuBmiZBPQGM3iiN+Gh9UBM2a2hb8euwjWLnUJxy8pmQn
xXwNgHW2JqrT8VKNOPyYeAVQ4R/FSRHvjIwj2GDOxcuS5M8jHGH/XVDvS4185jLYAZvHL1LeNsey
wQ+DfCv9UFWoUIktgoBFyEh1ph3zGRoASkLzZvf7F+e9TFOggBGjb3tXvcHvn3JC6c9b6V3kVHHE
ywLwIhycthQAf6TkgzU10/1RQBz7caUGsdxiBaoMAugFKEbcS7szY0GvSsED8WcZWQVDqEOBZf7x
YO54dazVwJdAInjiL9R5m3w1l42RfBHxq9yxOm/L/SMO3+4XSDMqJlECrhhp2O0allJ59wcEmPhq
8VjfYkG5ZuadkTlplsIjn6/s1CXn8hN6C9xDkYqOetKL4RM/iXXvED0OFIcPEe3lFg/lDoP/fTWO
8NmikIpfUbLoq/vrX7d7u+OdjzbIf0heFx8r3qzXIzPl2ENA3mj/HlJvswsa9aX18d+gh/8wkeJQ
o64+yFGH8/pM3Iqy7/H1XkmNr5BJpJHQjiDp1pbMhjbzZMti48r65yT7FSJ5ZfaLaI0JW94guD74
TPrb8uaF6Fyhem8DSIc1+9m6x8um2L9eQqnKISADSOwB6vk7oxw05s3AveLvDTLPO+0bR7hfvjcP
YP4YNQ9m3n+6xXEKXAChGeHikLd4BlDmQmGrZJzDcwvkjqKPqDG/H5vIfh5/jLkZ/iasEHw5XqxV
qLKyM9xdXlZUO3O5AtU1+fbMZ5dA/szXfN5yBvY5P4YmBihtMeHmfTYlO6kCOLYjopaFRtg/f4Rm
uXi0AUddr9v1qhYTBBJJ2Eo7JzvSx/kzX7N4Y8J7uD8GJ0gIJ+JBbBDDz6oKdeizWWda2c4GXHXR
ly7hLpahKnqapW0X9UmFlvV3M7CIazm/UO33zkDQHh4GVHtluoiUAQLVNrbweZoNdhg8iwBRLez1
SuYf9qLiq47VO65W0luMPjwvsNVRZb2ia39bi78LMhbk2veLYVli553UMgSr0ITHD4gK88ggBFmg
CIMB+OoAV16FE10n6TNPslopqIQWy+F+doHowmw+l20JUzwhSs1dxP8RrX179aC4GpT3iKY6OnTA
nZIHoNsSHfD5Nv/gvMyynvWi2u1bb25iPKf8GHkhPuqjJHzM69JTvD2Z6vPhJ0APu9efpbp1A/QQ
eN3GMHbFFmxCO9+U3vF/YfbzHJBkJpMPyXy0HvkGmiC84mIpS/Emfznq1tlfDEGXYb7kQHBWyfS8
qze7XD3bG9MvuN+9mV5xnQ/tjyq1jhnPFL0RZx+go1PXAf2qpwsCK3Yhl5h+r4+QKosl0gPugffG
HPukML72StpTCb1jGaYun+nTYGRvgf10fYeOqHbI95SZyVw6+Xs0zNUBPhRSwacFDczVnplsMHK8
BT2gkYsQfFxoYNnT35DMWapR/WNGKo5mEsHA0OJzkp6hRpA0yFkzjkmQvqst2EC/9t1CVqv6cldR
h8yMEkof9d3HZC0m6GaNUSszFaXE06fD3Wd14Q9tHAih0mVCaCbVt7IyaEv816S7OHUUNzqLGfon
cUtlsdCrYarzQV7TNOMvt5O7jHhtkNty7DQlTD7MuQU236IH9bUGh9oPuVe6lBW33HZEX8B65c3A
Gqluq1Nd7QOmNf4Hb8qXjGkvUVkPiFPcmgF5nu4QQTAjC9Hvp2dx5QuHNEfNsLLD5izn5Kfo/OAL
0e8veZsJqKyDRoyyJwZ19LdJ8HIzDJarEg3zgMOPcsp6jkoWRzlnOUDHQfsqbDh0CJM+Kjyexozy
m9WyexT4ipGZEx3N2RKzTj3+lkz0YDApDHQbvxu0HHUh8TOtGb3zZdKdJSF1rl2CSI7nFgYEk2F2
M+93DpTWzAovH8m1sV652Mi45/8Pt5AKYg5G8DCzwUNwUyXLIvtTB7udAV+3qFq9E1PWb469k+ZR
elSpKyW0Gx7891B3NZ4C5DC33LSAhhVQh5V1QECr3Fd/jjeVB/m+dLwf76dPeKBKFp5d6XAE+gf7
TY0C+mtQQmXKxIXRiMacfUuYPhYVh/kaTCEwHOrWDTakA4+VeLNf87f1Zy3H25LMiNG568Z3psJH
1zgdYI3r3SIV/p06GnrIULHL84o3JMicaNuOlO0pPh0ZD+nL8gFGw4G1iRVKaAq0H64yQFjfz8OA
fJ5MhQqGYUiJJO1XCUpuhlQokm2vhgUFgN3SozmAfN0+uUk61rj1paeycibfcMz1+6C3uxuum5C9
zAIFJCtHhPO6fTjoh55EyIZMKWUmIfvZk7H2xsraNyy/mfSeaOUE0l6YEf8JrHIGU+kbXyj52Emk
wUIMuMfbf0IJIgZglp+8CxbWwkurmKzahqu3NGBqyXysTR/OkTWBDVX6N6SF8FJCoSbEt7T5HASg
qtycrCaTw05dQZBvh8zNLZp3YOLfN+AVGefomsGs6xFT+ArJD386Ad6iZKFEITrCo6ugWdof082M
O5Birhh1cKgccbOGt+OQtazZJQDtp4Hnu0XO+1YtpNjOQDQ1Q2lch7bYdpCb38x7uOYv9eS1mC0Q
pIhMrTMDrsNxfghWoJx0c39ITfEpOT4NV5V6Nb5NpGVsqlQG2Tis5rSYN5G2Fwx7Xrk7VzCvw/RC
/8SS9AGmwiy+8CLHwYiZ3R3md088WrniRXKyS23IdcUrmy/GTum3cn7QF7xNJvOuNFu2Bf0pugkX
bVTZntVND4s9We4f/YEpyfxCRRs7hJ95SP0AAtJBwo8GmBeC9+U/pOit3XzCdg8SuFB3is3o3/R1
ryOkRMls2sbnktP7pEzX6HpOThnV5wnFWDEUWVYWZx0LFyMerVWLc+HFkVQugvOla+SPfBse9b+D
F/UGDguh+5yq8uN1b2b/VOysMiHNreCdzm9UkmdJdb1atnFjxksY5SUuZ/tVS505e2GTt4XDIb41
6GyRQsGzI3UXvIfBGonHZEqhAdqVE4bhzgi48ynGYrOhETEpIWkatovPQGOUCoY8HWwRWUybnIwn
7AS87l1ZwmL4ljboN/htgDAiDvkuqSBtvvliNQe6Q8I1FoWsfPYUppSendOzLm0TEkl0dDkJWn88
jux/o7rNMApvZPNOM9MxGyDNCm0/DeygzlwytryYWYOHFf86pVR1rVGRvzvRCgkN8mqdo6P03oBy
YkLm8OiqlxQCPL+P+ttWw9VhGRDuUixYCTVzViecOg8J2MyBd9vz6ifowIYFWjUJYVl3Acq5JbdZ
YjwEkJPlnvUQ26aVwo7mKCW3z77Zu/MwAZ9iyNRJbX1mzXDVdMzHsn5kN0QLzRyKsujelKFEZu47
9G9U4s9Fd78XGB/Eb2uIP6SrC+mkgeL7mLX9bRZNElz0Bs9saGkU5kKW+/H/urPbtu0uB5bB0+CR
+Jf/ouuIeWRbGi7hg91uedTYelecwZrRXvZfJYR/AnrxrAZgR80WdnoJZcl3tuPL7Le8NWDWUA8Y
kMbBP5sI+iOUX4+vcobLRvgU3HLwUSch0bzHR+vMS77RCPhhwobz7Ksj3i36iEqwyOT/5g9nouQS
FQT+fiyoBWwldC2nV8JjQs4+ctizroa2Dzjxs2FWixUTvsIjcrtlOPAQGH7Rh20MRQi0osv1ReOA
/Ujc3pBTSSUVGet1uBC5Tk6919Tg/yq4lQXDrsbUiQLY2Yz+14wDcg3Ob8wgcalwEvFqfqn4T5W1
u16mZHg2viCuJAQO5mZGOR5Rd7Uc5EZ1EgN1qrIzSbbm90Ce1K7lLHR8TpRglJwSouyJt9uXEe0l
7bD7GGkNSayWIErzcSvEs+CsXD5iDK7rBZrIjwcL7waWixJNI4QHKZMqVQAhzivMHQCs1tQliEQL
EM46JL7EKnBv2Y5s7IFFKfCdd4EcJ25ZcldMUsqWYe9OBhP7rd+2i0Fo/uHR/S2ilQRzp2tIJz/S
Q2geBsqL4871FF2whBRz68qLZfSibgqBPsZ2VGQL+/KHKFAL9f4AKFIdU9320ujz+ZUwJTXEMfCP
K0EO9mApsc5qgFtwr+IxzCK6V2TZHpdtWZE+5YwCEcpU10Yk1cNeSvQHaRUeCKQTYgcgipP11lA+
T2t7lFBrb69mQW2d74I7meK3qZQCEtTYG/v+RYtSrF+PbDlfzTpxGT77t87F4ONsnH0Xh9/DzUl3
VMa4Kk8ysOa+9Ei2tvEHOCXfQXRgKjmjBkOxsjwF28Z+xW5Wj4ssvKsUniA7V9c9Bsc/lJ3zkmQc
cyxuesxgbCHx9RQB7TSeosM+cSRmWsQ3/HSVHT9pwSM2nNOwH9vBDFo8yPdsCzAEgESW+Q81f98W
Bx2t6Pxm3Az/J0rFZ5Zcs0ZgqyxZCvI+yC2HYIRA8Csgm8aoibdU+x2FZN2aKoQ8VAtrfbt2TmGc
PFUIOx3yqPDT4FH6+IAbUfuZFSmbaDCW346FENnZF9J7S8fs4ruH29HAFNYy76uRTayaI6ufWSCg
vScnGT+tsn1ci3tJnkmaU1Bsv20fzetP8SielaV1OhtzuSRN8PkTQgYvxla/XnpgfQ0tfEv1RqoG
+fTrWcAtaQGt6XuoZusEhlxlQUvFBCOC+8r2V5W3G6u0uXefiEmJo678B+eEgFMYgJIG7DpfpWDt
mBq7FRMVMBy4avwv3wrX5cWobSFVQA04oIFffgXswU4uyzH9vwv/Mn+IzffRUCp2WOuynlCwRt6G
2np7ujsLbo8cVxyFYiJkiHVQ3xiPmk0MXKSCp4LbkHNcnZl5qNA7MT+6yCgEI4ZHHSuxpplSuGFK
CSZ/5ObTMSOFMSkL2CEGg/D1M58O+cKaVN5SoArnFQ1Ms1U/ASMyslIUdn51+1QemNIqvFd7iSk0
5po4idaSZeq/YCL0oIJeVkNmTv7B/RUD2XzZvQDknyNHl93YERzRDOvHUhtkTSHwpTi8l7RXmbfa
aIBRiLNRRkaP1+5SDo83YrzH+J0dksDT2q9tktg+lFaVhI97DMoKG2/f6M2/dtixflx19vmYUK20
Kmzz162aDO77OFgFFWpZ7PI+ie6+dvVjPQ0lXfVT3G0t/CdAvj8d6WxTAXgEuuGi10mhqkDKjeRl
LCQOqQPLoazqIkC3QkrwTqPsBTlop2CiPCa+4XQnl4K7H2oznjNz3073nNtW6Z5snqcZtAXusDee
YIB0ItenDpuwgcsJdwB14xTrLitC7twLZJkS/rC2Cxx74sfvv61pRDDTZikks6Ho9IAB8wknxHlU
kMGOOTGWupP09eNtA5I4crA0biqus1yNVP0LLrCGVw70MEdVcELHjGsMh0+SY9vZD/Hv4HNO61Dh
aZz9cbld+sITnrbGaC23DzQil5kXfiVTXPH1tm2umKZ/EPtKtiBfkA7iw02/bxoE0Q7X6us1VRDq
uQt1ESm50wB5h28ZQav3DhxyQuTqVfbVkPyIuMVeKM6bGsiqEwDFdWDDbdvZkii2PVtPENUDmZgG
3colAUtgR6MUgA+dfJCf4oaUE9li30afGeaD119zHFMbrbfjVl4FCLWcRW5zALccW20U17ZmSzcG
R3ow89wZnwBv0kJ6ccdmxTYCrhiWhJqeuksbIuuU/LE/dXwL3dEOvpTLEu+ROag+zRy5CwUIx1lx
2yJWgmQ/1WnnSmv+T/7WEEXV7aAbGdIxIDWwdNHbhHBmIdsy/4nO7rb3rqpukvgQQK+eXaVWZQlT
FChlP2go4fip4FIolhVSGGq06ELKiEz0gFc10I/SI2bQ+iQRsdCA+/3vmI3mAyKyVkZjCsHe8Opb
6Z3RBUhWgNjThn8+Jqjf0JJBhP38QPm3Vn9rBTozwCMgIKa9Au7XAa65QFfsn2+49ytxav0+GGTb
Z0tzM4tq4tgdSx3WRF8ZRJ3xCjlY1ltd0v10D3gnbsNwCp1FKIPTf2Q0dnRBO7aB4FwlnYZH3E9u
Q1Kkd5KZZIgGcWZxBNz+U+QrLvP0zuex1QFUpz+DEqJhwTyYrBJEByj9cAWw3CR2Qg84nmVmU5kJ
QiBQHK52U/2/x0gE31uAuaNDoUOl+evH1EjXLeQqV69FsM36AQfLtqMXtcu6mvZariWC6OsrlewS
KQrdbTU+G8P27dyNb3ExUqFJFMmBZa60wex2pGr6xrALk4jif4f546T14HrAxTLh2sHJPLv357G3
XvAjqypcg4PqIMnfvn8qEe3Bq94+JYNqffQ19bSXhl7BAYbJ+xNkUR/ofmtf3A1fCbV/gf/EM82W
aklPmn9t/3GMiNTmjafq316hBA6BMOs/8mV8CuUMzrIHz90qCI6WMTI2s3FtTT8/F8MWFlHBNZHq
51JjljDDmBLLfk0/G2k/hOMYkYNrPUuWgHSUSht779YS8kiBIExIK8n3o0O1I1uYlqmGcFSPWqBj
RiO5DB1Gabk+7XlT4UrawBRDVjeiwANkiDmsAa+9x1G3I5aFx+1cgnJyzNR690Rx0mGTEfT7Cfp8
/SlkQ+CW97hu6q588AzQCaURCiHqvIsfTBqQoVt8vrzCpssCyVykx8Lk9hXkqkZaACXkKoRud3Ey
WGQVu9foxdXbi3Tmjy2HGp+D/9Q3z0cFIrOnIJus00XfZtXOP+sG0PwIPaJhbhKW94zPmtB7ARXK
D9Bl5gJ8tQ61oUswe1Oy1iCsBDdTZl8Joi3avkRuzmD9KUWvFaIPZUD7Mo0SIRwReIONZfzj9OMl
zsjSOLwsmxjmR2S4WcGsMlFm1q7Na3Ke9MIz0P87YzdZP3POWGypyr/pfg2KwTyL7OnFoYM6XfSF
7ZMFoYpc4CE/hVw5sCncvjV6Z/nZEd57dWzKoYf7tAw0HIY6dWoVDvV+bAIQBvdY7OAUyHwBUf96
H2pt/KP5q6V1Wjuc20V6kDSOTEkdEsp/CZ24i3pnNxwQgKtRJUfYwiKuP3JZY/J4sHvtJQNwowti
LFygB3QoPpiaasVooF2T4zhJst4WygM0+HsHLiUnZxjBsQa1t+QT+T/As9YyPi/ToEDkg/BTJiSk
Vv12tZpL/IHwcAOLxfmRk/CjomfCYAf3qCkfzVcxqzV9mt1J+we3qKZbhBMnydmaV/UJeCX5NKYI
HQd68pnBWQsNW1Y1fbfglfewaJXmp/PGUyhkqrFcCBRzBkpQAx08DiaBIr2i9zo2cQY5xCe3cY5A
I+gFu8CoUn+zgR5/rqU405sr8TQW81IMj2+V7c8jqs8DpWG4Dy16lWn/W7YqFtoX6ynkR4KJpiR9
9X0kI9YS9raKzpBN/Ojp3V1t/qCYALbNqElBe1MyLEjvvAzrF4dzfZ26G7ijI6Cry8gWnnzUiBGm
X/JLsDKV2t1dVHBQJSg2tRLFCKrr1cw6UVoeYiq5YBlKyp00N27pcZIq9tewJKZ6nXHoZ2LekWKB
qatx94zItxdGdnRveCgecSwOmFqiyB7ThnnSw8NgrXbgaKB7kiswfPoN/y7NcaKN2xhwhjytTlCY
QpNw5vABzhug9CBQHU7mUNz09I2TPYU+zE7t8pgpTJZRA0OuvlCedKUG7czbfI+2EZduYnLYrgQj
VipL/0MfNArj0l5j9bG4X0roBa/vUhYnGqFV6TBSoXIRy+sLdNL9ieFyhhJVWQRsZIYV1SrPDwPv
wRkZ6Bwz4EmZZdRaJwH5P6Tib8Q9DmOhiDUkdT1+p9k1L4+Q1mJmIKHH2Qe/9RQF41h632wzLNOc
pIAS01ZfyQVccrFzOZ4qLnSbx0IGCN0Owrz6WyQ0Q/cjkBFlXEzOU7QmvtQSs96JJlbXcwNovCHV
9vRAFOT1BR9rp2h0FFZuLXwYDy/Oxm44q8KSHQ/etqDuGDoZUYjU9lnWIHnlJCPd6GlygBUJXEQn
c2z524+8shIRFUYYLd0Dh9R8xrv98BfZsDbxLcr4VWKDMTjDVCe/MFXVb6t6P5wMFE//iOXvWquE
bYXwYdSio0jNxTlQRXaGxt+bpN1MTTmA0NeJNrs3db/SKG2+/JK5+D25Qe+X2ERlrYL9kWw4v+Fr
1QkcBUy3Ao+rmI2IfbyZUYCcJGxVg6u2tTScOo8s8EMskkHqYJGgiLpBwoFFnzRFYsUr1luLfBsZ
jQ6YRRniNxglAhfXGNKoNap3mtWCDc+eaufp/NxmCliuo8aM3OzZXLfS2PZHkQoxrBjfuGWKCmJr
tLgFYxeXcY1iKB1UpNWz+SbGgenVbc01xvtB6MBawPm4J7YJktInzkKzlGKKRpiNGjMEPz3zRQe2
JeuvIyYh2BjSq9R3sAePheUAn8iJ76/PlBLE7BI3zXPpLuteVN6SWlQ0Qep6pAwjM+Vgpxc0edCl
wW3S8k0fDsxIvU0c9+O8QpjzhAdX99BIgMVDE84PYYsu9xag2TSPg7sQOeGaqRXT/C2PESfX/DGI
6Gp8rvg03CN695PZXjV1oTu7KHBIvdZe63UrzjYTM/6lV2BhKDxrR03I5LD3pu4mQQcWMd79t2Bj
brzXAxmi2UiEkn27hCngpx2jBB3mbncOLg4ixAhBNax9+qfwb9KZEtp7W64JAT6zM46NzANcV4f6
bpY2ETlzbq0n0dOz99gG1FJXLyRs3m32gh6/b9S4kMnTa6GqsTWAYJUCTz7LaBlS4WKNYuFTArdS
eFpblfUGsA/0CFE9gROup4voEQqRt4kemegBzI0r+M578Z0HsBK1tAAvv1nB8y2RV211V5Q6toav
8KXA+T5/1HU6bh9/VXPbCVB9y1G+JFvrTXdB8ptah7TyHAdI35cAF1L2wPrysILNx12NlXCFum5J
fXE9pmezGPDPdZkHKzqEMQvYer8yUqH6xZYrHsLUAmaIyc4FKEcaujhoyOCMXkceN0xXlT/4kSE4
1RW2iPYov15Y7B7CGxywzQycAIAf7LyHZ/9vyzKmgA5f/7ypBdkKwk7WkZQmw9B9TM2aV9P9l+eY
zcEn4Z6resdW83yZBFLAabOznWGe0dm6WB19yWX8r1bxSczSXXClhq5SDxA3zDOMldbewnupvwBP
CNgJMIRP11cYNubbPw467gUgTFrSkl64y764aiei485oOtEg/MMuE5vPyXG/BKUlQe0GZQ1vHWvH
FtlHtjsFfcVLHLjUw3GSWd6RtKw6H2GxaLf0iS7WsZ2QN1v2BIgTYyl4bfC2dL8jOZmDjL/dxSE8
KlQuDaSC83Rn24NXbvwGlNZ0be0WRVHI0PkfIkcIWKxiaWGJfi4TRtSmLsoW/WBcBk/DZ6HX4i/E
w+JTRBePqQrIiyuZA3XPCZk2NgvyTgQAnuRtKUlUXGK5bAzBHWh9KIrau2BO63pzGdEUT3P4PNmr
PesTy4OLqqYhPLykIrzDFEJTnOnPexZ0/ub9V2lt9zYc1cU8WiwRi+hchR1c7QU7sm+ZGETWOH4v
x8hQuWPKwDyY/v3XxeZuINyhEae2VKdDN/xMKBlFBoBXzdmopi7bnx/4YOr1gpskZxEFycSkqNfC
mgGXua4vmTwX8IvaZh2kNkDsnwcIzSqcs6KhdDp4+Fqk3fjW5lZAPw/jQJn50cnLDqahG3qTV9CP
3m2xOGy+cPpICgALbtFQyWAyoRkXzuOiFfwBo6WBexOg9KiyLgEuKYg0g84DuvbHPjwRWhRfGh8d
wn+rdPPqCcaEe3+5ERvh8+nLcBOLY0A5llP3ESiqvSPEL51ge+dhpv7Cs/zFB8vPIsWUDkmJ1D4S
e1QOdboj3P3IK7fz0JhZnDyXXwWjWsSvZs3O927455TYQLYYYgTMG4Fa7POpOFcg7Z9JPBFsZlNR
p/o0XCHWuHxfMHyQcb3A1CuR79/ElCD8iS6q4/7cJ52ADH1wEQU7IpNjid3IIygwf/sbIbcj9ddw
XRc5xOTUhHipbmTpR9BIu1WiLU7dBsc3DXvmnipkE9w/SuHJay3sz/1SQaSEG2m7cez5vK7mlaT7
hltGzTckmKpDf2Y0w3cKkKkyAVrahdHM2Ic+8paQ9lMMoTfyoo2v5FdVj6Ojy4dz1eM4dS7nGICl
xUloVVcaIYGVMlJkef2ejq9YDNytRH1lXDRp8K3UDfSnUkXM1koyGnvwUVgaE1LxMw6u0O/g1q/d
3b9Z7sBP6/GrEHMkYA7ytqomkWZsVNaQy7d2MX7F6jd90cHnnV9KTsiwP4/D+fOv+Foxg2KhrGeW
1846vHCE5JZnsfo94PQGrcb0lzeXs/t1Qml/H2fZAhoVtNQaz/kPQRpkTCtyjjJvMUzjV8NnYzr/
enTSIOyuUcSZ6PuLCm9yAfdfuayPOPJMygwRJxXACiH9sp1cB4KHwuSbBLzZye17+zPU3VfYY+xi
JOE22+IEcV7+uFaLwOD1nwYCGDxbg14LaTTaM0rXXwORjM/gAnb84F7gpg+g40MfoQiSxTmkDJiS
TMi9SOH237eaLjXyo/c8sOWklJtcTNvTgmlhO2lOoglCd5sbbV4UNUYh/Ga8Gry7jX3CmGH5qrvS
0yYu/S/RA0g9jORsvAuCQHqd7XndpVsmlsM9Pd2hiGO4PW4T28MDPaaaEjBAomQrS4tF29GN2dly
hkzlbHevqzUiWyY1/BOObwt4R5tB8CvQy0kpLo6o8cOK1hddCp2/Cvuzz+NlK4ZQgakiqbpl4eoU
7ESJWX9WEgSADetmextcZ9fkabVV7D0Y22AdL0Cj7/h7fNnajKlxTUh1460HsxI8qxIPXsByAtkY
EEDjIxpTS4G34yYnmveR7Bk9X7roW5oU78I3+Ct6oz6cf9nnjd+x30LwlviJpEqRCTgmxIN16M1I
u54s4VhM648w0G7gYguL394GxGcM9ezj/0tSDo9q49nhWdZKNN+ij+nfMtIGwHURM+5ElmXn7hsw
/5eKPKHWX6r9ZKt8d6W1Mvzm1BelIiLWZYw+nnNqrzblailTtlZFPaY9eL1wbyJzByok6HLy27wW
/99iHKMH2pbg8oOp4TjzvQyWkpIP5ra0s39uU1Jt1Fq8iBHHOC6W2Wd/jQLOFwMsCsmA8gdFuhwa
itKp0rlw7480EB9yfHvWK43pn9fnK+bFpquFbRt/Esgnk32IJc0bfGCriNHsLzZB3sSjprzaWPk8
BWgjq7DnSMILnsOqxpmxMtO++RyaNoymJCK9bALCDPzOwNvnc8xJLLOxh5/citxniieaaZ8EyCQQ
cFdNkIh5wZju7Ol5vpM2F1q7/lCw60wRVj1VtExw0Lbc/5faMDrO02Eihn53nzN5ECSWBey+dg3X
IrTcF+elrBZWv/Td+UPjEhQ7bVcZhWoNyT94ieOBP1Yr11O198tDkms2cWY4wdcShzASc9lctpGM
FS3yVk6DqN5cRDrY3mDfZvYey5MSoj8XrGZLcjfImFiUDaNZzxlmoUUdXkamhBRE7ANthFUksqsV
yNFBf7Kv2ip2XG7fjeJRcpeOBZC4+gclnPueX3tG6RsMqdV9PLd044TbiOn9s/UdZlEWXBdA46Hj
Hh8YE6p7IwlEYYhzqqQpH/ZbfVOlervh8FVSqja3D79yNPbd/2IG9E8HfR31qpMdr2z2S2mFoyt1
k7xeMgB5czoHgGnQvX6ZQL5IS8K+CDMG9pmwmC3OWIiT7//a6OrXFLer9MqFwKB8fXbeAks0IIMV
+NyoglxY7w6zXNWdjjC6TvcdXfwzXi2iER6L/rGc28gTMzOhO1V5T6xZ7YUpRiF6cha8uZxRbKN8
zp2zGnQ5GyQMuWdWEpIWjPaMCgzHj4FBk8F6hs34gFfV6vH9TkgaSeiyb+vGXVvPlQiYT3vRnfvg
yyvptgqdnj2zbB+Wwl1Cf9Jxdy8aWyjjPHITkdpTOdljLx9Zr9A2co2NnWQnPMxCdVYR5MG7Q6T/
FvS0oCIoS2oXG98slRGx5ujJ5vrwZO2mgp0hY5RrbWbnQ1V3PWASSXMxvt1hGkuA9q76gdSlkdCs
WK9sJ1g4gNdqJMkD6T4MJbSqaYIQ6RerQZxV1fgmkhxMnuDHmpo6YAVfRvhQ6uDZ9zvrKvwKo/mj
gruw1q6AcAzk0nKSflkGbvov5+CFXP51nn1vkATszR7ufZl9A0b+DTL0Kuj7gJb8I4r/+7i94hT/
3cMyzHXFbXxqdtrNzylEDLUKaDNjtThsi28OJHMq1MO4M8OniNjLG3FCzak7XfmWWV03kZgVsuvV
bhvmSQ6DsMhW1AD/sT87uGoWzcU1qa1AgpsJ0A9LnA6eOCm2FsYg0XFCMN5XsMe7OlIxsedh+6bJ
R+A65rabo3WESwQ4UQ1POOthJgh2O/QkSU7bNS5HAxU9z9/PLee5z+cu6m/feFPc4FWvgzhPoyJZ
nyWUgHtqj71QC7vEmkwvcMXA5v/1shp++g5FLDPiJd8R6ojOjNgNac/dSOgjh7T/+X7EkAh7r3Qc
nv2eEP0A7aCyuFK6LdAGhqzEs0HJKwj7o1PY3bnbNWHYNH7c6zKqd+5uswLlBXcL6H6bUR3S6Qhs
qiGfkuoKCuTN2tliFFhF0Ir/qVWLKWXUq+6RLN73HhUYtBBgGkAzF3UyPb8nvzjJu1zGyZOCwD3+
wbag/KR6bBQcDK9mJOJX5VSQ4IV4uyHn4CXZnQsGu3BW/2aVDuF/5nhguq+4yOQUnIsgfNNr5Vp7
9yxdr8H1FqYvzsZeuDC0o6Bwp7Yg3M+nmGoXWHrcc2TdxwyPVwNVmGYEgcVVKJY9w0hcWcNcPQME
0KEsfNmqCZxW73N0+nDGR3CmjxnACEexb+f23znz151O59tsEMgg0ZxkHvWEJnDnq4ltmnepz2ea
6YCXNgx+V0ueX+FE5zQzGm3ZoeTYe4AfyECAioDqu8EGqUHLUxQWLJPaZBGy+H1rk3zYXaTlTbR1
+HmkvWI4GDWBrvFyNaO5PYLjndbVX0liI5SLWDyAza4D75wTVIGBzrjnQCarEp1IblskYl5K6MhY
PnkRK7WD0AVF08WSvveCYTID55tbo0to/5LgnoWgvhNCZAnWjbBB6ANY5ccFAsPq8y9a2igTC6AW
gsg5Vv83ixdpv19aCGPyIZ9rg3K060sJM4+sE3cKUk6yM+4Tc8XfwlLV5reSGhriBhPqCa2OGQ6N
gXsUWDy9Yfs9N8hcyhFSxcvydGQLdqgZLM+jZF4EH3qnUTyQqCNQjVBN5i6ii+ReabkFkjJ40B7T
MwDnCRh3rFS73wS4jzdQpTWvjgKYBmqqrib8zs+c7YpJHnHQTT8pfTQD07kjvAsLbfQCCTredC+k
smSyoWmHRgzMfhWBwtSMAuYQTBxpUhUnh6bp+LwSYzO5h+4OjbgD08tvYt1LdKupPW0AehYoymZ1
vW+DN7ogVhDr46ru7nLzXfNql/S0z7egrj6OmDFJ7rqtocgkTBmvBKmnblRNvjMgREbGojhIcsyJ
ChSX3MfLQnKk0H/GbTezJB3weNxnYxuFQDPPKCWBTwnPmvq+a0jMJmOCj+FMPfgi6r+CSLi+Esho
0m2vOP3impxybOE0DOF2Q9fxtUvA89kXyAiyz1hQmwDeD6u+q9e+5zrbnxIYeXJC76MlEATwlx07
3VX1lFskwxc5dBgJTHJtOVo2BbAdCM1+8gqw7O4l6XUf8XOWqe6PxIMZlLDW2B4N3ngGX2fA/X+G
t5t4B+wIp02BmdAX0xtBd1sBtMlmHRb1kea9izWXYKzQyzYhEXudHLWp73/syAvHS579zcPY0x5D
e6U+zhK/aTRA28Q5SQEffyydS1pSdAPDZXbobT/xhUHBKlfeki0Px7JNqWaPNMFIj05EY+VEP/hx
n2zGoS0pB1VRvtxFkZQ5SepXPBOX0T9c6u0qTqzLbKdT+NCIDfv3Oi+hFCByXS2JyuNFHQaTQPhK
Upor5rCbI5zc1tBcvEwy7RFBBRDX/6NGWRLWgBIu37F2XkhoEfQ1mtBZVFVIpPRGrkJPVdNWJfR5
GFO/YqVIAGFpqnJf/s485QnlPlARqfegt1WR1eVSk2jYs/sRczo0Z9kVe9MBFYiC98/LIkX05SLc
lvHRoYOZmdaiAapPSml7PaDo5xUjI/buiEhAl9dPn2lUtaCYfR5JOUaHDdbKylSjyX7tf6rhpoul
K3YtObCk4eSytBpHIlPJ73w8mIZx8cVk6nfKCwXJaCq6yKzsYh6y3QpyQkMbuRL8CbhS3A695uu3
UTi9QBLY6Uz/o0b8MyDGKi0kZshjnrEyCH4zPu8oWAvrIEIdit/L0hKmuft/YagTQ81+jAjBq++C
arFiGEVm7r5rjZQ7HMuZOMmkNN/dJVJqXt5PEJrqRHyMeIOQU9Bg3bBS4FsYXA1edphh0Oh2l2oF
nf2C/TsKNjo2nmvHJJAtl7Zhq+Y6zy8galt+nzWxocN0ZL+mkztPSaGLGpz11QgwKcvxn932Y2r7
Osb+1Mepd4Cws/LS2Oe5K7zDDlucj+TMx1YksShIQtF+MzLZm2vFEg7q2KeV8ttnvppQHXLLoZbi
Bw2L6hGvjF0g8uoC3w6Gv1gJktt0ZsDRRYwaqWkt/WldeHbqwNxzsmJnUdq4xu7lR9d8nPqHOdTc
r16Ta+OenjzO1IqjHQiLVuAfUio7VWevcq+mzZ09p9HVie6us4RZND+ja2rE2dReWe6npYEamHMT
2S0vAbW1BSAFBHY7JZQ7k4B0NCTB5+60pk7SPvDItmMfQ1duz0NCw1wezHPQekKjQ+4mJ6HB2FLh
raLpFxRPBQoiWa5E2iQLOhUH4+D6S+Ihsp6+Cqu30r01Coe8u/7hRBhlEBCWuMFoYCJ01xz7oiy+
UBdLA+MOr0/jnw1Hj1doJ4fBczCtaqbyHjmBan8HaHzXxCV3uVUspFlnfjNgljwOiiFzhp90FtbF
WOH55Gm13NBpjZwh1MNyS7M517JpI4v44I2lCA0Ah972vJ78b265riDpgvEXGGlnJVma4WbHgrlB
/HISEtuQmm5psL25mERdxiPcRQQ+aBWuPn9sTW0HGDU6L4IJXNq++PX0clSzfLZOkjHmF123WC71
GolyUP8YnjibBk6Vn3g4XEeIC26r8an+Wp7qxw9luacSH2OqIqK488GxaQ1jyYurhsaCpei/rh3I
0sXhjtrp602uDN4wAlSBcJ6mxN9tVpgZ7e+fo3xUQGO0HN48S9qkuyYdY1X8yGucBqIdHap2ia2x
M3tRg4m7szHwncGzs909zUPl+gnOZhXH1gt/CIQBWp5nE4e3uZQYHlT/WYslN7e8vCoLkjxvt3YW
koj/VJUu2kERUTVVZzgCJbd4IM9kncOL7mxY9yYIEC1EG3xkL1p4IZ/tNbViN0Qr0soOvpEZBLAD
TbvOBIYImGBW/vdtwz37FZfZELc8/ksahpTrrxXv0K9XazpkQFvgvasNNe0SaYmQRRgd+vlYfu4k
oXeAfcQzUkNkBDxBZpvAUCpcGUemkr3rW3igj1WWbfcZTT0otydEMktzdHElzOC+pCnHuuO2zjkH
VnbFSuvrwE1+Xuau3NMyXLsrgmI/z2Qc1Ubz5vbaidmiNWprMquhNcRfIV36XI5xVA2avRLVVj/4
HZuSLqhvWk8wjIDHWf9Y48i4e8NPkb6Qfa4yoQVY2AezT4l9kl/TwY0W7zbyTG4ZUvKtrOZ4gRI3
zmGIHN72TP00VIYeRKc7Nc2XJsDZ3Y5kIhZXF4gtSMdmvPYBa3xJoenQPkxRWp5VL2OttAIQxdZb
KVbta7AsLrji80tWKxyX06gehRDyiDH79BjPluqxtKuTDuK8oAwlld3K2q3mYy6lP+NHwP+VC17b
pAuBbGtayljAvKnt/Aa7Kj9Qk5HVyYPIagXDA4xir5KoNgwUldGY8NMzkLTcRYuV7K5rNHA9A3Un
7AFQsNvhEsah3XgfYopGfX7f/f1CUueWg/Kq4BWXJRO+6XzDkY19C7SdIQRwCip+O1ob3gdYxdmX
mxr1o/jiL+KjC6Ymw5hE0PuVlLs0pefZpJkYp+0f8Q/sUwVnbPy6NO/KXZ5BSaCcF0U4RTVOe+zW
w0LCV5B7N3K8puPcRC93C0sY7hvlUIUOez7pJ6Udd1OatT5vnRaaB6jMeivsT1YC8yxiXmKD+5iz
FmoeYhDM4oFB5ASpKHbVFJKkBNiDr6iiGTRdh3DnN9oxpzdYz7Uv286gZ25KplSFerJ40gSll6Ms
bE7ezTP+7F0NZxYaJ2/OhTvb5UUsLHkc5XpGO7PSZPE36a9UWAmbYAO5Jd7zhuxfYfm24H01AOmh
gJQpOIZYDJJgFnmIh/BzlmL8pdda3D8IKpEhZM/oCzsvK2zRR3yGoKxBCydWkkxOQFpib9EEyfJj
VPgliuXkW3YZOg+HnVgrMQ2FMTa6HEDptRj8Cq3//g+sqBE/r46DMbssyqxO2OjnNmjWwLnMSGO+
pr1OXA6HetnXenUumg8BwOtQXGg/FwQ9er5itsCfR8bUBIsMgi13zb1csdvF7r+ppUVN5EklxRKy
+JZz/LT4COWMhlKmzxAGfsQvTjzNoQf5WecIReD/7In81LloDerqYsDOlrbUUMrMJNf4NLFfsmM5
7g1L6YaFBnX66Xg9PW6rOwSvtlbxkaoKZazWbsLfkBVISvjDMDkXJdut3/G++ofjc+WLDY0W/XPJ
Kv1zx56eUmU5tLXrFBYplLKIfl5eoPdx5eoB+SnfQTXt11xvEHfa0HWCc+6YTQaf1h71CamocYwi
oIPY/20IBXelKt8Nr8+9+IXq/m85+ZcSAs3RFtVWxO9y+gV15SsLMiS9pr8sdeXtQ6LWJzxT4lUX
RnL+JPxtiPelVbt7aXU5AAv3xKduITFq0A1I42j/ygez/99hoin3KPKdwb2nZdJl4HOi4/5COnSg
DdXfcbFJkc7QaFqm3UUUFkZv2a+sL1nLEbMsFJs+d4sGnI+y0VcM3P559Tl2+i1vC7wN4voldir6
Hx+NMzjdy4IaY92Qhuns1qwlkvEApGizkrXeh7okjyyb6iajaFCi3GhBIrnOJq4hT/z6qraOb+mD
oHSHBNsZ0oaVLUrL981fjCnbT2B/lGZ3w8V3QgzhfbKSrOj2jesgqcOS/0lcx8pfoPRa5unUq0CF
iY1up+B5J7mtReXNQE78Hg0JdnYWdieTPFKpgRKQ8HVKrQ8asDbcueTi9qlzy85roH6nAE0UtY7o
16eLGOa3mAWyMTjcSWBel6fUpqVTppk3zdqZ9N9Ltv+rcDu8sWFKxH7AwopDqISFxsTZDgdBzh9q
P+DO2HnTVRcXBDQamd5LQY2UJ/aX3iecW0AGam8A91J0VMS1nDQyKWM5J226T1dZagS/rr1vu6RU
uCso5kDZUJ8xJDg12I2/x5hcJItpZBQ8t8Oevf38LrTWYB8+yhnighws9j4V2ieTuHPhb/n/c0qG
nRuDa9APnw/JDCFxxtPNaKo88dwiuZIptBka0wNUmXuns55qaEZKcutje25ZeLfcMa55T1am5Q+3
KxeTU0g1hfuWpr7pu+joDJukz78gwdekuS+LuqmFve+CNdXGtAggU9HFVtKPl55jFHMMtCtmKS+m
eZVywrQQje0Cq3uT+ZXcIk3Ex1vCGkCX6tEkFwFB6l4iF3w9mYub9+H9dkNPxAXqbcu35hMeEEVM
VdqyWoSFRTLdjfDiizD2CVa+iAkG2DjZ6udp0kHDp8Nu1RRkkG14gyilEGoZcc6NcxnDHUHKJeV3
dGwi6IBYHgbBsIEs/TA/RhqVY8npph+bdHfjj3Hq7TTGuRyyfMqjERHhcYR8iGCAZ1VW6puYKPYn
A97i4OrMpf3cBDZ2y0FQstb6IUISn3vwWMFpCgVwvZFVSJO5joJ5lCSL+7fjTGAm5w/Pve+QV+wR
g7r74BIo1imH7mXG64ebB8iKD1aUUs7zYlRCDvCLhVOwch1TwQn3XRNdyj1WB+AsPnBE733vhcSB
URrK7UgTMeWfPRrRcVVsZB+cOW9G9jgPpqK5gSfy8YgQsuEclCgadtONwvEz691w/NZmhOaYU5yw
IvwkXnCSrMXktg1KadK+y1NcR7kLnsTxhPDfaH5NtCHFD0o60CRKOBxJ3WHeO9DpL67UA61/uGE3
SdhlM74PKvAHqhecRLJBxk8skcIhWIzWXq/VWhuyimQqvQC2k9c7zV2I4hPkC3Z6bJGcF0AXTfKl
isXYoxkyicJgJBtswuQteG+E9TvzlDou2YLID4tiEMsPZxg8etyRJvdcZe11b1OhawrjSjPF8omR
iVO3060LtEFXkrY0SFY7mVgYTaDVNPOh2TyhSF1u0N1r7tlVfFm3anhDX+MNTvpLO0/8yTbr7jPZ
WcxPZjyLZ4IHZQvVn+IF0qmsPUFGVVHVkwPo258vzQNJbjYIYe4uOn87TPFFVZsebhMYZt2SSM/s
3/e3VBTV/coZsm6rWaaEP2fKeDuq8zkqdqMmJlHVFVXNN3JjatupuIcJ2ZWs0Gji0X94HjGq1+rt
S8vYixARaD7BUJMWfoCWa4xbhwKhqxAONa0jr1dZF4XEoMhIWoMrVl4T7kcOWSLhGT6kyYxNHktj
40DHSFGnbdyjU6zZ3ao5RWtAI1VB9bYa7fQAUGyQf5beMhdiTeD55Gr8/xdAW58rP2XYBHHXtlqt
KLrMYeXzVHnRwEnFJSMtPdcp0WCaJ4GMG3xUTVr/eCXkUTjwUdNErir4zI3s9p+92PPi93KzR5S9
dJVreodnCPBL3drvK0Ve0ItRupyTWgO6eTkDrun6/Ys9aTRvaHxNoEP1ITC1CIGWd4MhDYnY5+18
Ph56OOTiM3YjKKsBJWtxigVcVq71Am0rDZwG2/gz4TxY4Kjgy92stc6nYPsfWtx0YMVeC/ZMed4X
BJKwTTHldOR2ue3/SVYpCq8uhyREULLpKGCM8tNSophCEdkZTkiYzeTmuxbnxBUCLSITTat+G+gJ
GVk1vjrlbJjq6Hz939tiltyxrcZzPvsIIusH3v/DFqqgBrWYsndoVZLuLlXm33fgubPrQ3yrIZAi
yKMzva5/bfvkjK8wkA79qylvs3wllpOVINstOhafyJTPxjllQqJ7G/3Mc/GUiM3Oq/EdHSSm1uZJ
t5Y0eM1JneTbK+icelsgU1qplUh0zXeIC0ltJHdhlDC3OAj+BBcV9iJC4HX7tg/DJszdcwJPEgrt
xHqC3i9Gdl9uyqCiUEDw7slmiyG7fsEjrzaaVQ5Mng98/iA7Uha55rGUoto9NwxcHwL+4SvGKKB/
tO/A8e4HZ0I+/USnkJJtBjGuVQB1Fq12o3HU9J4Pp9Fa5BEYQlqon+U1gE6v4aECvo2qO3xllh3z
59Je1DmNKVEQLB4xctiRRlTk2y9Zom4+90sie1aEhNbup9oPczvQqLIWt95kStzkaHWDDNVLXCNW
A1rxSgGc6TGnTOtWHQ7F/CPM31ho1SITPLhSxDP0WzH2Kg70FMMl9JnwYeKZaGsVHjmlUTEGQ95N
Ax0yT6DSJoBo4nRl3vZgJ9EN0nBgMCsDCbpaQOrDC3HDT/UVXbf0bfl6p4Zf8J2+igVUx2EZu9ZV
aOwvKaNfTYYveLCa6ibFae6YvCRszkvZy1gNoiFJRSLD8T6Rbbv6jADPQHwWy17M85r/jE1gStU+
tVqfjlDzxB+mk6iRElUuUC5wZK2KdcYGNeIacGz0m3+6qDVHwWNzgs4jHEHIwQcdb3USMBhSSs0l
+CFXJTP1yL+cOJjbegrKkmfvHLIYC/GK7ClbjJKyTyod7TO1IH6+bpDDyiJLBGt+SkYZvEKWJoJQ
p6QvoiDlJbf2OK6KmXCyw0jw6CHoekJC9f+98lBMvLeXznkyQJg4TiJTs3xX8L0nhi7aooPxbVM7
jlrQK8jH4bN5UIobxolbqNwqnjOy2vcD0YnW4gd/AeIHXTDdSGOVTWwkGESeU1Fn+4JMskej8Hcz
n4zP9DcGFkpjHYt+ou9vtbRvcCpZtJFXQ8+x4OqFitoYL5msQRc5shUVpyA0IbfIzWBfz1yZa4wn
WatYl2aR7xnwpZDBwOWnn02NJWaRv7Y3u+Y9ufji3B+dor6lVasvluIESyIgOw9Va6Bhs4mUvjdT
/li7zRVw6oTjnRwMyu7VCBZYrjvgUnmjjGXz/h3m2hRtHj2256vgZHmlM2FX03HnfJt+uCO/bNQM
EUVaHLrtSo8ISAbrbEad7dt8M0jnj1+ifr5rINQ8TOrNehWZF1tCWrMqez3w2YNnZLMEm8oVVSfm
ZiRNpL+BhUatQ2s25pQ7NJVMsONBJR/NX+Js0HV2l5QlQcV0booqb70kdxDzZc52HNQFalYhBJf7
AVLakkHFKC0GYpLhqHFK7un2eTqyjyWUevbiSv+D2ePGA43UCgWrfHWX1AGRaGuLuMdKGqLPpEwb
5dcxqVg16bgDv4wk5NvmHi+5/0anozn8EA1a+VOv6B4PrtE80qTb7NTumR0OvkYZeQ6vk1soD5AA
9pmu3r4fUTq1t6KPR2/a6vYRUdZ5tfWGcILnmp5DHycbzS/ZyAXhx2fX+DT4eg2vOvVZfs/Z2lre
4+GpMUNORbgYJC1vNaHsQ7UyeIAyV1pYAYuz4sJpnTjFcA8cKs9CjeIWvxkmw2rLXafttfhWeASD
nv6TCtBT3bDAmFNDsoqOd5zIRVj2+MaM5DRKLXhbaUONndfJXZgNS4PyNG3sko9gg28yC2sBLoSd
vRJCnlV0lgQ8Mt7y5uLvMCGxE5A8kTtvh1/5vU6I1fbvuAOzFBysqBC8BXm/qkAkZaUEUR8CTx1N
vu63EqUeQCPpY1DbZa+U3rZ0veeOJBbHiDwaA1Rgr6FgPeJKZU7wsKdMtTi+qkZ1Olg3D/rhjpwf
F6vumMvQj5oIbSE2Vwdau2sL8rdZmjEmnjf+4y6HrA4szYvjmnPBXn3pove+CZvHnuxDezkfnzQV
W6IxLo/Gea/FR4KcI4Oe3lZvsdn9CZ/qKJvHstvpM4AofvgzMbI6iilat+hl9u4JQj52aZvuzfnj
IqNsGHOVsapPCOSgdmYbgQy6lIiyv8YM99ahtxcj1X6CQtMfMRoVGX+bNMsIzCCGPrQGBqf4BRHO
tAfDSkLD/g2S9DwiQSbzTRv4BYzdRqhTOpy82Ofz1JEWsYmUzxhlk3OYYhTXOO90ifBu8KXiY4UH
dNDmPH0aMD8dqnQnmxTYxiYsr4/uHxGwbUhICOWHGB1K1nsMm181lMYh4YYbuuSqt2M8cXC0xbhk
vshKEf7JK+BIySvNAysqKnM1N/Vtc/9Qlhjr6HT1F9MVLSbbjb7MNF5uuH5IDudS9TV451dOLrg1
KN2ItFAuYEr8WqX5Dj1xPJDnEF+RY1jS8j8NqrHrQbIRUiJAIfGg0+fuqjggmy42gSp9JuUmGTDJ
xKXD+yb/Gfy1VSD9oqJaojX/9KZvGWjySs0hisjUJEgGsqlDl+DPoHQPhY09muN91FVx53XtSD+T
dlNHrdiEkdykDtJdxh//KFb7uv0LjbTkpdtllBr7dfSxu4PKXuebzjRzkkkbkK4r0/NShDDhgrsl
tvduFmBUeOPtHLmkoFXwtm4xlClvMDlTRW9r8VGmyxS4R1+od9gv+BwQUyXUpTC1rth0kk3k4Ts2
YmKx7AVOj+ACumN9mOKgkSOfiKxf3G2fhhiCKRVQ5h2Ni5wnoLPTeOEV6IIYiETx85mB+3z2LpfE
+t8QsQEHmS9zkB/7NZ7CHnoL9cRWTPwk2B27E9akoehp5yxKAX4uIdNEcyviDGdOw0x4Mc+rwuVQ
lSbr74Ok3PHVEQa8GecRjN6/psHunJqekUWLFmCYfgd13RVekfpD+ciuUmQoX7d86dVVrnFxdFhg
nm0FAuZEC1cf5lgniuz6AXAETUoZpVSPxAj6GEYUKK5+vmj7I57tEn1VX4Jt16RIzOsMqMpFV5Sm
UNqL4tfkr88fJo14Y4FWpX+WrX3MioUopLq8cr5O5ZjQbretou1p9f0ktCmAbinOSHqq7uhzUuxa
U9Py9oIGvvgVxxjS8Cj3Ou3jAh+bqufdKWhkrNfMcC+I64p66Qgu3Ri4V4i3JS+tGdh9IPdUSk9i
KfNd+O28vwfh5zjv6F/0mb3MnReNgdp+LpZO52nFOpzrAeoyaThg9k94vMILBLxk50jHwnOvG4Zt
HFIcljLS25Eu3Q2Cl55JmdHW2k6uR2xXd9mz9cu1MgyvP6IylCZOrOMCUiuW1wFJvCvV7L4milbh
rMpo9wZu9Y02AimvvZYkri9e9Ee/l0j8VTAu92V1+uCQb4MsPcIfKCT4xhc/KgA/p/2y/I0Iquum
ZIJ4mxpqxam38taQS8IlpaIm6hVEBI5eXaDh+/mND+fFHLGNrqcZ+hE9yFzMIgc7uq7UVM54DJJO
3OdVaYL0QBl7rL94aF0mPrmDhA+AILD4vSJZWZIRa/NsCDN5jcH6vRa8ftTcI3OfK5zQn5iYT4LV
qg9xwe9tX9WHkMKOsy73EAuZKZIJxEEfHMoDUl6c8ljwTJ7oBTv4wlmJ/Ev57QzFMs4d3y57ETnk
xSQ/zPkkLb79m2phEeecoZ7Qsq/KloeevpUxGb2DG2KyKGNIiS8IljKZDC+UrD6ngENAi0nShomG
vhxQY8bPqLtmGvzpfuHwkDR5nrWCTf26SC18ybIUyysGaEjB/unTHYYYH2Y31E6DJOz46ljVYE4/
AeOd8ndRhFX2RcmQtpieecLh3cObhu9Plt4mOvkIabQSYt24QR2tgtz6lzGPyly12LZuPDxvFf0o
1Ot77OOo50pF+CPCz+gwduw6ap8ANv16haUOXuOJYUccCKklI/4wrOyw1hrhGmlFp8Y9/l4KFAzt
6QjAN5a3/Yr865OC6xrWjX9LbXjbf0/JUzZbmEv/fCCNjLBvF2LASwts0Vw4WHiowLD0V8dsaelm
TGoaJC3sj2BUgQHVcE90NUUDkRjyw8LvRcSJdzlgw5Y1sP/p9cuSb/2idw5nGkfHQ9KssukdCXSJ
Rf3FM8kZMVszxIMgyHGrfZicx220uIdbFketlFGvM2c0XZT5zUTw0sTHeLHtKf3AZEZwWPjGqdIA
NI80HngaNxK2FKkmSi7BXpf6pVGYBQ+0NtznvGxT6fTlumBvidDfTI3BAuCjtU0xHPt8zrsl+mS/
WBuUmDC80jyFAyG1mSaoAlzfcbDvgfJJButthPnDn3BP+rqjUyzxBrh5V+AqKED7mNoTyt5KcLFH
KEdqvFpuwDOELEs7d+08tSnu5CzV4UuYvraIIHD/3MOfWTVsjyUj0TO0jZDRBEKy7Y5LBbiPaQ1E
3J663qzyzoUsi2Rp6o0DHjNFCcXlR1Iror6ELgUBHEYm65twSq6LNY3h2P+xKsrsy4j3ZfLjTL2Z
zGGCctxppnPV+RHUf7WlINbFoN6BlDpMcJG3yXAR3VsHJN+P+ENM6DdAOnvYo+u3DUMBS2h+Mn2/
Tbs+i0EZfk5rak6xCEt+whfUyhYYnhilYRtkHpTbhPZTwkt+pbtwhx7hLZ2E9Vb+hqfh39rvD+A9
9ykI2v82Yl2Er0VwoLYDmKCo+X6u2iJV/EH4Jc2YfmRW1D0DWUWxV2h/UCfPnuRBH+pfAsDtRV5W
DOeGiwviqy49aKunyVz/joDmbzJa55wnez++fvpzOqlB1wZGlADEa/mgRi8Mx5g0EkPJda91dC5j
kS4+nEOaHszZOk9ZpwZQEJxzSiWOHED7LId4Z5UFSxb5gNrme5LCn6yTPqnOck0/4exko1kj9JIT
+1kaIR3gFGwbcVkm8Oo2j/yGcsBum+AXllOE+THs3tRLi7iP34dCXyFgsk3v0c3kKFn4L+ztZ0uq
OPMl6vHHqCdICkm4H/8nCQc2KsGvDmcWITK6CB7DsKXb3ZH7e/EUisB0tTkUiqVzWVsM8CMdE9so
FCHh/TS7gzOlkIiT5WUJJyEYdS4LDO7Omh3gFs6pglZnhQEkWHvrmiYzgLU/gYR3t9TVd8QnU4fV
nZ8MjpcTuqP4UGMIA0qgymauwJTd/VrqTuYvDt0t3DbUfpna2p6+/s8aM7ZEYCag3QV112U/t7lo
EVK8BpCCQlxwPDZo+L/BtSVbFTm5rBYpc71fPuNLS8NG+uVso0DvRTHkfZVWf03UNvteCIVrtO/P
WFS4IsiNX5AYKkAsmNb0usUgjKdqwtm+bkxxOiO3Drw7BNswRfYBl4zs1VlWfgpLVDkTeH1T+Lqm
AcVFJX6pYPqYztzbUYx1VSuAIvwYZjiEynr7uDnEA54SGsNEOhRC4Uqn4Mh7acgTbKI4nyx78MPw
jA8nxMPSf0V+HXUR1V55Vn339TSmVICIxSXcMS253g7P8LzSyerTq4BDgiw3LzHvyuN8FNMjy0xC
dhj8GAGhGC5/CPhO+SHyi9vr+ZIK+CtsVZkmPxwMwTN+WT5tcttiDfAb7/vffkcaImUr+oemY+wM
uhmXYW9QGyqxiLI1UTLsNbTTWncrdFn9H8YIQ0o2kIsjEPXDxbC7DPyH1df2Nfo5uf4kVcISdleE
indtI/dDkCl/8dhLMQiFbiwmnJIjXvlGctGtGF//aCIqhpDw2YT+2FRwZGozWLpqYkU4EP1qluWE
ThwwT0krGWNbakMPpqu/c9DWzzDzNI1S6SjCoBbnEPMEqUAvor3hRDFesj3OKSllc6EkcOyVNwSu
3v1/OdN6zjoNhrybrNnIp77hkWUKrNr8UdDqmWRjS6jY0QeheyY3+Hsjl0yegx0xIS8wMNmKhYtn
VdIwJwQnuImxJhSbVbdmGDM8DzYJzMhNAOWNzMEkv+qvLYMdI3Sg5iDz5O7gF0yv8Fu91YSZoobw
Pehsg2pSOzdSDTVl3LCkn222A5Bbj+WOt9LHNb3CXH8YIacfFyD6IAaMagItBNQ6eZc7//LHvDK9
vjjaWmWpZ4qzID67P7L1y37wu5LHU1eAKKqaMUGyyMaDA37tGfoq15tZD/F2jzTQftPvPVSKLHTY
QG+WU0fTXZtONbU6f4ybsycfz855Vtzl6QGueMdilbmDKhPyf0r+BRRSWxVaApmPB98aK8u5ypZW
vsyPBkDPmQZE553rZaf3V2r9JYa6LiozET7Iqu+rmFFTClHnwoeNzm8IpI+LpLNxv9a9We/wbehd
4nGvCNvns8D8CkLrNvZrFBqof8YPYLMyIch20U3Oe+czyHO7HvzhStVsdeXfqPCcb/KBWQldM8DA
qOFunyYcNLbM7ePaK9OoDz89l2GVAy+t7cZJam/qZE0KQ0BBX4LTBNGKI7gIHJ30VrXkGe3LaFmz
GHPTOnzjUDJlBeBRsTlIU6b4C8CcfTTE1pN/5oPYnxzctY/PHxi00yB5V2XZBSlTfb9QxdCgXLdJ
tOwYWVAe1SZaW8M/j5GdOr89Bt0a9lKiyDB7QNhV34z1Kz0+loJies4o0CGncg+TVnte4rtC8F5M
KlnHcyFBejIFXCjs6wMFE00MIU+Cb8JCikEMmi8kxL49icozlyNx74lch6gQkkMrWEHIByZVvyvr
ri/aVA3wkEyrB4e9hX/ceyXvNmAA5ZLZVYB3kEMVL+cOul2Dsety8nYEcQfLQDq/zwGUk/1tuIXh
muzI2jP3eLc3nwWuF8Z7HVZUNzMJh48wXPBE+eDkyZYubHS4wED2OlmM2/q9BlPzG1VPyKx7ECN1
A54jg/vrv4y2rEwGhmSduuJGLty0uWEbwDAi9KoRcm02ZesaYjaUGPCkHuEqOdezT8DpCmxBODcb
sED2h4LOjShU0VhLBHD8GTqV8WVrkyIyX5D6GxW89FlPOsGso9FjtUQHKCMFa0GgdExldsRBjl9K
KOfFxRi79KMXyadYkjlis8qMNLoYcHi3b0g/gdOE/GGQABnkRUvzmokrqO3rZxcw9tvwXUXOo2rr
od7kTvWbtnacJoTFtPtgt2bQDtLzbLn1Q0HgQgs68eSAUnhunB7cBQot68EFRKA8DhkdqZ7SZYOV
wk7ZPM2jcwJLS8spLfL8kFklDLWaqXPS3PTJ32s4XO2CvInw3U9iRfCHKvTsk0cZstqJvxvOmJIm
jdwcl7Qc2Z3Au4D2UXdIHMZUZxkznkr0qb5oU1xxEnXYgBDNEHQBjqOV4nrwYDAhVd0BGkijezdV
b9idfAk3bR7jI+6jDLKy9nsUY59CZXpMBqOlXh29k4I71yP7DImvKnwrDm0q2NcZSXAP6v6cNZD+
cUX5W3kcS3vpUFQlsNO5IM76+2AeEFBBPDJdJqOcBjFqzALPZE4M0I15BVGMVJvEAQ6Fez4xT6L2
0ONgUHwb9N8/pX/+MfoWOmDRMWtsE/0hQ4gvTuQHFKqGGOW6HmdGJzw0UcqhFZIQ+AtZM4qDF9xF
cslUF3GTFOV+5UQYubulLC0XhX/FfpjEPWNUCR+vbnkJQGyNh+XjnIfy95VQOIQVrv79Fp3p8Uep
T6cEyIPH5WZgxrdc4PAZs/DSGUWUXumqvJxdR0cPfqYE00LbIfL0kHpZk8S9Mtn3j7gZFkt4NVsW
5dzB85WzqLVeDbApRaN/AAsNNJV7S6AjxD9RmSp6uTDPJtwt9MauUwPtuFR7pOF/u79sz6JEYGJp
bVOaS6Br5HQzWrSLybb6wCkre5HQvQ4uks681AdufargYiIrrX0TpAv12FwgaaGNXTOzL9zYL6RJ
fcHuTUcYtjQZ4IaDNBeFSN6/OjLeOCGDO8vpKRIca1o1+sETp+jdQbFcf/yi3D93NJYfgTJCFX7p
PwUqHQxRS6lA3Ty0GYYNBfPUeyrseqc9OeGp6FoGVg25D2VEOHtoLkJwlGnT3QrDjRr6B+jRpgH6
6qaiRRgf4dvyzMQPXvRLR63sXtNHHTBhis1ZQ4P08IsGiIg+mGUg1caWHTvq9gaR5OLoQBJFvXYk
ggwUx5q1BY+cHAz3cLoLwjM77rtvUbl+cxRlKOjovlw5z8fxeBc6IhoxVkrJ2mHrCe1It3KOZvE2
iVMa8St82lUGPHVjtySrgTCNczGc9S53VsWVc+URvRB8Z8dJWWENx/YfDP9pEFdCuz59P0b5u+Qf
w7YH2a3V6r4ZiX5hJeT/SbYKDry3BGqVUIA06ir7ig6fqAi97bIk+Rg8U/xsBqv1tCk+rNVplj8c
lQ+4L0f7q3sa0+IyH/C7Hvjfw+fOk1SJiBrJz2HtyLls7XLukGSDPKbMIZ8FVkDm75xjboPfNMom
di0sHPbj2S7VimY/hUsoDrJYsPGk9180UxqL8+Ki8ALmpOVZfrNDvptGsZJj+UHIxaRPn5xVObDy
nSGkQVF89DvrJ+VL/ZYTZd2quZr3SR+D253EC2x1pRNo522fJN2e6nUsnFGx+ghUN+d9lVMyIXaB
YG4tLgJrlJP4DLXWQbKHzL+22cqHQzgBH7ej/h9ims5z1Xfqha7QniSS1tSGEENstsq+7mC1IgoY
57uQ5zQ/QePQ9UxLQ50Qm3RwFD2E/UbPNHXZ1RFRGtIv/DZXd8/GW4YdgZo7TpSNg0C7PYed4cwT
Fcv6E7I7cJlGTBipm9AMNm7tYH4gJWAXcTecHNnm1M7HgbtCPewaPakb5OOqm/dvlubd1joajywC
gDkDvDlkNfMry4MEHXCd7JyQ5OrMsvbXmpnuergbc0ZnmB1PkJfHQ604vQbN3Rb/TMBRHEMxj/oz
yRZAJ70DSdfdOWZ9Kl4Mionay/f9u5MoQe1lGVgqVKrfEYSE/YXfSRyhX6gZpt46QDz+DP/Xwog4
GXHXuA+a++Luj5sI0MQbz7CLI8dF+T6QlN8ecrq9deOM0q6TMqwTUIFrrR7/h6+CbquzbQ/ZQk7M
mMBE8+qx9UGoojMdzE0PGopysTyF/k6Cm7cJi0eH74dXjpA6xpUho6bFH3CyBce/o+dLNMIODiQh
Gq0w3CKLnI5YMTtHvSOOuhQI4RiDX6IolQO+lgFjiNj3xO7iaWALBraG7M+k+5piLGjWmLu625UU
0w4c2VgtmBMHc8WS//O5qMyft8k5fteB9ETGb1FItfXFo0CPunh/fXLxV+O/DWFMaDF/vi3rDptG
Kqs/GwFgng48KzUkT5iGDRnsI64o7PFuisomMpABfPZQtXC3xX35xog0IkgDXpFN3roDjdDTeOLE
9BGU7eaiwsc+ClUnTqWqfoKm2bxiL5jZr6Nv1uHE9nKzKCHffLr++eRPQlWp9R4iN6/NFspIr29R
Lh/o4pxPFwZhzAXXDsbgtKU0LIJPb8KxBAuswrSwK61RiMARLYtCeFuGmx04bdwb66jS+/uEINNx
GvX1U9QO9ZEyL0l4KnFap37+T7LlnQACYBA1iiawtwEse43DKDXK//7waP0vlK6NFzYhlX1m24Lr
44G+edhvuEx9rVf3X3YaWoa+69AXwiXQaylkq66CHdmYaClygUbf9MbGnOKtkrTD7zE44RZRCtvi
Esqs4v4aNVfc1pmV+LMEzvU7sv+n2U7EHG2hWX2D4R21dMKVw9OYkYDNb5PtHG8CXU8dskT3yWLm
fgzjS7bsrOL02xM1HFQxa6+YR4fj7uCCibz2BuwuzNqHl4jCmMuhQzlDiAa4g02PeYM1tePkTpOK
X/AtDyYKIVC9ecAR4cQmub6rm11pwR0QFnZdTwTzgjW1FjCRJvmtuM1wScqSd6gzlTnuPtspmND5
nHFAhth97cJoOk9/Xi3z+sEwJOdW6qRIkwxEGQFuRYa3ae6ggoKWaXBkSjlvxO9XjQB3QCBzE6lT
l4x6izblhWwFBP4F4SqiM7OqGSBOxWK4LIKd+IB5fTT5jk7siqre4eCHAi7+hHnIMooUzN9OQrn5
X9vSy+i9i27x2XstQbOsYJ83+BAcpXxFzDPo23ZIschumgLbMdSocyqPBwv1eYkyaY9On3QCFYnm
M9uhGHLqe9A4IF4Z85J60kIkBAawr/rHabYXzMQPIpdWeoCz5nPkqsgAfrdmpltn4rmQiX3bKFiU
MS0tOof0zq3zQqKvL7zN3+k2n2T1JXrUlQKM6n5mgA2ExhNxI6jRqADhvugE0qsUz5GDvotp2Opa
0RjihmQ7Ai77/gpxOaUIVieDkpmrI59FZCrvpBEzlTloY8SiT3/b1xZYh7dPTC4pqFZQk7GYWd0g
1FxwNaD8Wm8lR28uaY8ze3p4oLoJRaS+whoI19Y7IESgzm3cBE5OmS8zvW/EwuuM8TRNxUTF50W6
EDYZ5fPOz+yy0U5mJN0TmB+a3wNuFFUX0NGdpglcqLIKJffn88FiU7UpSRPXxNa3IoYK9dM1uu7W
U1pixfOFhtk1IZhyavUiJXYQeIGGUfyhORTg+yspG9A4SXT+clz9De8yIakkKN52Y7PPgVOeAPU+
+NSKPoKw5VAVxj+nJ+DxcKgCZixrDh6K7nXuPezr9FWCDz5idlYAWpk+aUufOkAZyfxC7tARWoF/
c/e9EHpPDIT808Q2Na11DREzJPTxeMAqfEYmBhMgkhu/AeteHeSuNlVnuO1T+w0tRBzv7Ult07qz
crKygR74u4rqs/1lbwMRZoTX2LjsJ2J5fkaYt9orqwwDgmcYR7C5n0biSqH5HdsAIDHub4lrOtwa
FGM1Xdnav3EuMIBD9AoLRVPjF9IwOf6czxuDnkMxVzkDsgciy+UlS1Jmvuj/m1o+mVS2oafwvBob
W1eUROr3SCKwpgwxY6+TxltWg8kn8IFxLTx3Bk4m2fG4YqtB+DCxddCjzkCjqNzdZo1lMziku3Ma
9yj/eGZvz9d1KPm6SyPgXDJhd5VLHyUm4VnO1LUdpMVqiE3pR1BxZFvWVlTU67PMOf1dDWDLDKTz
gxjBl4uAuB/ZoQdxipox8uGYHu234Nx7ZQcRF1J4cDMfZKFmNxm5O5avDnCRZE1dBlMgRYbhIw1K
Scrzfewogd7s646WKBzuvGn+MYhp1LP0Ecuo4mWZmnDiFS12mTyv+Ppp5EGV8vfdgAO5qA3QAr6o
LSMHdfjj1qazsLcnSDJSn5vYkuKeqAcTMVbEFVMp1npV+6g7XxEBdQ/bNpmeASGYBYeKopSbjyCL
IYPD1mB1/iC6wJLE4V/ik5Lz1RP+5umDzHp0mgArJoT/kgMNLxH6DwkrOKCf4O1mVnZZEsbAfBPx
Dyct0LtW05TqMjTl6vhNcRBko5wmlFdqLvKQde6nNBVMCVWXj7rNifN+vJ1m5UuSgWIOeGFXiA+M
1UocvA6fJFf1MEZEE01LVilPEWDFvLiD/PJ9j3CgUMw2h/GRUzkvwgsoSYkY7+xbLfbchsm7zrZb
YqBhHU2g3vhaWJSOJ5eOn7JQzAIbry6v56lODUp3NSA5GO7PuMTdyxIucfE9iW0J17pkxlOagRON
JOp9JikG+1BPLGmHtw/w5kWMwGsRjED73PSUg0+n66kLf3t7WupTQ5huSHJuYs82WyO3u8P1TQUT
/1RJsNYAGMMYwF5J3xYhw9Oy3lzEcF7Q+GGZgCLXHgLAFju31an1duieBEsZUQhbf0C1P0UJDmvz
AElqrqPOohJlmHoBuk4UmegOj2pwZ3lZ5RFS0mPAJyh9/gWRKkMR39jv8RTWrY9tVOluB/qTTRop
hbHHKwvWFqKzu5GpwrThcHFgmNshXasi+kLpD8LPfqNRQgpZi9YKyyBk6vrlQWHbSYo9+bz59wH8
yFp1GoylA19evSNECqggY7sJsJm3qCR3vYamUDnGQxO+oY6olQ6PAPrstqLciRSSgeLMkpYs9BY5
aTxqR7dwTYPaWRmz/xfq48Nbds0pzG/AFeIvTTTORTuus3Ok+wobo/t3aJmUbbWGuR5M5JhHyuN6
WXGX1tPOYISdtbCFdvSaanPVTq9izd60Mq+GmrI+mwqRlS26Qz3l+YFo2LMuRjFogPCMC2ZhECz+
TxgUZNGD6fwrEB2akHO5SDVeISx3OImFqhsbE9nbw1HytWiHkcxnHdH4W7TWOo0HT1PmhjAfrx+k
cHILMbpZzO9rEZSjD4gZfGwDMlZoTNgN6qQsHD3SuPQooc9yFXviN8homunAlz/u/Hvdy+pZoDG+
PEASg0uaHH1kCajJJjlglZGPp7kXSwqniFTDHX2Lrky1P6xbAS1cjUr24L3K9vToXFkml6jSp/dM
5hUVC390v7qvDFEidwBJsIzVjFMfOQcBU5NqjzPLI1o9YgpX2bGjuT22Z/nmSDeRdaVIPyHQNqDK
Luow8By1bUR7EmVdhyoKQ9Hc8VN/6KA5skEa85yyyH51kj8a3C3fBBgRg7oHry/vBVmj75xG0O7f
TnitZo2OsiAwPuNuoU/vMp1SoFG3Ska2kFyuY3G9n9+9liiU3At8dLWOkMIJJb1sil0LVOhEC2/d
nqS3m+RsHNzaQLbH/VNDnejmHBxYLywgCFSTulqzFILu17n7F4nh1FES/gIcTSeCtKWb0Sr1YU5x
CeZXKgOyLdWbcsTeSqkTLSeFAuBqWOKDVHN74v5ATO8JSC9v0711yeOd4Y0ciksKZ5Gx4xB9yIJL
dhvcrIqhaW65sH1cKIDzKvg638jk/Tmh/CdhJhKn2f4ot8Y92CTHGhxVWLPFYP0FYZXb3L15yIxO
KUSB8N6T5d9EU5ueOFFfL0QqTwNN1O9W3VzfLRPTlZ64KUAhGMLI1iyxKwVg4Re8qy08osXCI64p
XduV8IxwHgYbbStGywbzxw2/d2c7pnBF8AJdJrNlcKey3ZT0fFOG/K7566ToNskh62iXUvzPzrhS
hhoM2ZsDxldp8slJrXbnsO4aRBNcYKO9r4u7xG8iKh6CSt7NHzdhm3g4Qu6c/Wo51hH6m3DM3+xH
6vcU8lYRWOiEM7HocAe4iJb9I7IX31SnJ2MmeXSrpCxkKKCvVYtE+TXfNtIPhA5Q57ogqZruacmu
uUDhhtBNT7wPr+MpJ/imtgfr4Ldr9Fij8fXBqbUe/fmeajkgeyTt5u7r5k3k2zwZybQ5U6ZVjgAA
+K4Xu1RGPtGzpmbo4Bej0+lNzKLmfPeiZrGPL3CTvQbQGxU57qRVI8MpkqTsvN1DQW1momkl+nK/
2qwNOaObGSrPt7K9n06313D2iOns9QPwmH7OIsSLFhc+P/SWhH4uF5gi8WwD2Oh6EEr/TKlot44g
Bklt6OB6kJSZL6j+EwXc7qf19zcn1PqOAVfs9mcfI7UXXc809DVFbYQ4YikuHDBzUyRk8C//7MT4
wjq9mWcERab6bf43Pix/WskLQBdbb5H7Rvl1Dhcpp4sSb/LbzqxDp/WDUASuIezEGUKjLVFPS5XT
TRfhV018B5qM6G2Bqhq88gzjqwVi+6j9Gs6vpv3VEhIhXBUhMCkccP5Pii3kxK5mcsmHlESX3JIQ
jLxikab8ixPvdqKOTg4gf9UFhjso9yOeRlimbN9yoGrjTm0x80ybMAoQsecR+z1LsDKM/dWn1DHV
MGA52mP19tqxotpKYKeFPygc4SFHG8P9p2YjpVV6wrLxvV0PK5UAJ8L64lWEftKrgqFKKGbeL+5p
UQkbyFlLVmpX/2aCCnXOGn8JTI4q0plm0+uTrq3EPUPjRY9B2pw2bu7kyNFI1fsir3w4D/7b3sEN
rbnoUqecDenjd/rmrUJqX2hs/GGEhOSTvb0bAo9uUZB6a82KCouq0C+vXzo7IMKlh6vg8bDJcu6T
2CsrmdKfInreeyGi9VQNESqJ65pxPPmHGROLnjAmvVyvg6mMG/FOfTOZGJR0HsB842Jo+BL5MFlU
mYCTbsdmEEX0guGgK6RnPF6HsmiO6stpwruXxN9+4Gpo60r7KpbvMfA3I04cguvssfCOPCyDXlAe
Cz50zZADDLtl83xUThyDzxQ/Ike2X1H46aZL5TML7LhoLEwN4qGnlkuac6tFjk2barWc5mRo91PV
TuJ/JN5/pyHBWJE4ALdtKngrPfh9yH24F+dBLXS90oWjwyKZvRMvJ4WemXC/rM3ri3gGyfqU3ICJ
XNIIwtii9GMc3pozsAVBUVYrLNM9/pEJ2jJ7L0SnX9Hzi9pxfHdg+2lsr7I+7DHRDHMM1c+e/K0e
0vsjeUs15eUXhjxbrEfbnBBAkVKx/3j9zcW5JEr906Ic0IK6kYks22PLQqCPT7VdWqEZD14DTF1K
E+jYeT5l9Fg822uLglmeSynlXQYgEatG36sVOTlXLB3E2aHx3mpsM1njah9Gye67PuNK4H9l38zD
kIJWdH91CftCpbIlqbsDsgYzz2+fBn5OV9hVlsUKAzt01Wzv9EGbqQZ/xN5/V/1vsg3OkuYZj6Or
xKDcRSqbsoA2WtOcN2aDMeotMYwCti2n+kAGBxOBgj7y9NQUCvwTc1aOaTbyeC1/K77h9ByjpbTb
rECM1eV3brNMplC+z6asl1aVdepRD4OhmAITM6QrED8QQ/sxWYM5VKGAT91i6JMHOBwb4Iw3Un36
sUEZsxe3/MzTuHfXVEBEEBU7/WgLGLw8+FZqMkahpuJRlvoVREHwH4IJQRwR1rGdEvCg67e79Ne+
zY+blQ8+Hfbc5dEgKOhqzJ7imN4N12miX7K5rsx5N/Qu4VGD3yk3O72rHf2R58DEoSBKuKGuRkGV
Kwab2v3jR7JWsm/WQC4AVQMPhHZ7f5YAIEP0tJPfC7FOPiLM42Ombkrf6keXtISr1yRoE1c0ykbc
M4wuvPzPGMA0v+LlxldD0EJ6gsLHXTdf9J5nX86gVhNEfLAfGhYua/amnJXk1T4xzt4sFMo8rRoT
0FjasGcpTyO63HO35Flm1B7GecevkE7nHjkSA9TCAMqWpmX4JP/J3Ft1DRODmFLo7jNrzaM49SDW
MUrLVFv1QXhW5rnELRaS0HLRJZPW9a7ulex/f65K98aQHX6weZOdwKeDmBlyggLZz1+94dhKrQa1
BlpGzzKUIVnxPoFNJtwEhE4CQASfy3k+VTa0VH6X2I7/N4VO20HaaHWbw37l1oYa6YDjvg+4sSgz
WpcsRpMR6jsxkDuDPyzLE/8s/MvQipQ+pt1sKNf2ouAbB7yfOOCSR/rlPuUkZIrFh9r6EPV0BmB1
sxKNYUJr4VU3OeLWoIwdmjmftOmaBGY1i7XTy9X9cJn2em5qYVVpAXGURnvoBhHhge0e2ioIdgiH
o+FMt6vD9J+B89MowfTKZ5ujchnSPMyxGOCf8H73NDYawyZxNbXviLlcpqUNJtw83wgeCSRM0p4A
6CoOJYW995dimKF2MeRnzW68AbU1wBP3qKv2E1aQ29lMoP/qcGKG/yhdRXcrk5S3MXA4Pw+oI/lC
fcU2HVrrxt4mDyLqLtL5bsqRKX8NYKFNusO9bg4ec7nBc15Euujb11fXjIwDlswZuGDIBNxt5aCc
cgNNG+Z15v0uzBCW14YaqL0i1wUTZQiE09B3e/2ixCyH1mKsQAROUUU48AXWSYgziTEi7gOUBsH+
kWbJbwGkDn76rak4+N4Mp9SKkVqA0bRC2BriAAvL6KEwFeLZnQ+/NCFl86QUpjbGSaNdKP2oyaqG
QfcqoagtsXo5G83yTVfnXGIT+f4/YJRKafJQdOZdNakaB6sXseDo9jPVd4bLpCXdHi/Q6qMI9AP7
jX4/Rrdjd+4BGey5uow7D+4EHEgjSIOOT8K+MKA2uPBeHbLYB7nxJG7jY5ablh+gFuet9arIaDxx
9Xd0JDxYlF5uCZdUHBP9iaelBHebHCYtbpgPnf4KUU6Sw3Iqd0MxRNpjS4hRfBxwuHZQNKrGARVg
dJHr2H1fdz8n5YNrrhzYOcfIT8AYxPxRH7RhUVwxyofgIKNwEtwELA0yjoDzNTl+wDKzRA7/OhNE
pXZAZ51VaYOwoy9Co4eRinNviiKDOE50ySGCWDcLYpfCK9lg1wn9oJLLp49B49omEkWAOVh+gqRx
D9qDiAjOJnN7hiT0UwVJh3ElAvUvC73S3KefoUSwd6qxiDowNL20dgnDkR/8Zt5Q+yrlvZFnFg8t
qLrJgmXZAcg7zzd+p1H/sua394Mm3EIY1IbcPBZrXgqx+38rVpXQM8zdVjL3+GP/UTJcmsxc8Gyt
8SDdpHW1dlSN1SkbHFgQ9bXdn0R3EdnSO0VjRL+UIOJH9QKqldnHfQSujT6vGSArAoVP88tzOZv3
PfUOYesy1tySAW2fHGygWET0zwlq4fgF+z3qLrvlTeVrjTnpNGG+XYc6VRoyYNwiUGPam3v+fJvM
elkpU0u8jle/5KIN4LsFbHtH1W4xgD6ohJu2fHidWe2Rr3bD8G60FDdRF9cp1+9uafghq7zN+GPY
HL5YpHOyE2hjNzAQIdiSNDv1aGFvfWhDo453OSx68GC9iPBsg7X5+phnfa1PTK04qfK+T/mDDMhi
uGMxaZ6aOaOxNpDFIpGTqy+iHeQOJ8QzQMKI0Ddeab55wslkzDAAnj6lnpGkPMjj7DEbEDudFp1p
97TcRxtsry4bwmNvk/oegUCZu817vB5PuIB6zxQpe0Yej862gtzs/FJHZEXbKjLdSAF+d0kQV++x
7REDHp+cszMBtQ8G+X7EDvRzmVToHekK3VcYYgMNcv84DoxLTb5KRrxIis6iPsn+fHugAI9hCUIf
CgdPuP3Rq/ujb/ywc/CiDv4IzaQ3ZgUYRdCj/caa48Ov/0Jgp3iw7H8/a8zE+S+dND3dgdCeW6nH
GMvwegrZ2CpeLOflVf6z380YYEknXK/mmVBp0RcRgBVoesL+bZxlHb30FucL0jDifpDKcayl/ell
6q644KF0AMZx/WWNgQoi30Kx89HjvVMoAWvor+WKYQypUYMnF1HwKBO+L1Wa8A1NuM7UEYqzE0Wy
ptt1R7v0kodbzh7A69VXrOA5FTK/46Sola+XiJNx99DL29thW6O3YnS+i40JpoznDQILFr+qh1Fj
ULV5AKafTiE5XGm2AROgGeYQyVpuXwEzP8AMsCR69/aag/gk59wKcBH6gC7pZvVRyelhc/skUjLD
2I7aggegXP9o7BL2btCbT3LaAwaIeWtoEVYwnGl5QvQc/PioVCt6+POAkrBg+PmcuS99smxks/2L
3U82igtahGw0JrUZTcPgK8ObdGNT/wtRZpvjw75Jr+jmS0BjweTo+7fh1bGZCm7KlMdKyv+Q/TC2
T4DwiWUH+oMF6RjF2JrCqtt5fUFxennbikOqgXPlkyq3Jr9hXu1dB0PKQnEYry5vfKZEOVA/rOc6
ff3wtgyG5HNW7n/Q0obxjDLh3/+Nwmp+VcrVvJWW7uopddB+kNl/1I/9nVqMesKWt6XkkmoZP+S+
Pt5gt8/7nSUjbE99hmjraZPfERQp9zh+PhLGltKM/iw/vygPbtt8oTEKEi0OfIht0v7IQvNU34+6
qU95Wo26f7FQLNrT7N3HTrmwbApra9oGgx1wUjhrWnQObIevJpQAmXHM9ZADIH4esUasp/+idyFw
TiPox52SwHj9iLcNAMJ292bmCBzwHDP+5KpVc+hV9gYArww63svKuKvGTgCnnxsz/nZaFZjqwKWW
aO8qCJnmY0Bk3wr8LMHBYUwTBabzjj0XO8nOTI8BpSNFcnPU0lI8UNJFpKVnnHy0loYSSikmBtHc
IK4qJGngaggJ6+z2QNcQ5ryYQm4wXlfnFENVleoYjMkZI1nB8PK2ecL5M+DUpzz/WzSXRTyjFw+z
8po8JkySp6dBKk3ickNNXxcaTpGMSCkC9Bq0fjsNqQwY32OFPn7JkmoyHQQVEwvbT8ctdCElwOtr
G/WFeCLBfdXEWb69dyyAXZMR5AtR0Y4wqLm1/ilHG4FFU7FFlo//vHrPZjms00wTM/uhMQ5bcV3k
Vg/5uLX/HhCCgLUA7X76R63AGTMt/k6Lt8VCPLb/CSCePuuA8toj8dGG05tL30OpEQp3fk07BCze
tssVzFRjbFrNmyP1V1z0Njk4U3Tf1pMknThcjYCI6Q+ELT/c+gEHkH/MBWhX84kj4vC+sUzwXO2f
z9EgKYcaGs6zPaNCWDPACMal6xiRVPCceVve0c3NW687PkChHofmg7GGcgJQRSSwmQ3+GzFAUHRf
z428lXHXU8T3hPew1dAYDAMUxVz/zjVQ9A9Pdzs4sebWUB22Zls8a2QUrYoWHq9EtPLgWJp0GSm+
sz5mnCBKSvrxwxeTZfEhGt/xbC1NWPewK1tRPtzYU0iZg54dZlySVVpO5WWmyQ8P2YT9tVES4V8B
VS/hpY99jrbQoc4797Cb0mzwzm4UrXcNJNGsIx9aGUDMKWmj39eJFCvrq2PWqBniKDW4Lf1X7YaA
zsaA9kcJcKcY7suOUhUOWgFLcfdXPMo2ixoBl5sJZNHImahzzZH3JnmOV2kG0CE4gDEgqquZJeup
V0i3xhI+O5qUn2437eEvf3sXyndJ24xTVDFtWE9JgDgMUofPneudDJrtWd/E26BBCqeJjWtQM7jB
tYkF6zZzQM03iM+WGkF7sYr7tgAoEd52eh0hpop3nEkK3DM39+TkKhsXaJwdzPHzwhiLUYI75m9C
9jC7ozZaROTJkDKV5GFscEqCTGsKwoXQOYx13y64KlV5p2tzfmk3i9Lx4GsWxeTkbDkB/YsoiZMB
R68XGWuUSxf+UW3yDRHHSP/YZCTNrm66YYLucG/z9n/eJiSaA9JC3U3xJ7dXQjVaHL8SpjjWEhTP
8zi/GQwnb6r1h1rBoZp/4LSGhHcc2tXnflnSdQNduMrvCNVsRJ0o3lhSisdEUG+SlmNygM8PG+Cr
uoPov/lvYJbMRjkmv8qfBett7ANRdVdLxUiydhFhGZHQ58bFBFkfN2VHb3u49OrwXN/TlpLugDda
7uAUCNRegFzIqq2vFsuCVCfPwRMyIE1uXnCkPrg2S2opnsNgie0mz/0CmccM4Hk7qJvVQlv9bxgA
cOB5W9Eo732ykgJGXI+9+29l8JmTHCDyNr8m3eMDd5XaNB4EoLI/PgP04sD4CcRvW7Pj5x/pgC6W
BB7vh8YgsO8/p3DWElbrp4uzDW1SQLfRQt1pXb4+JVIRkEAt75NQZV/KFi7vgELISUejb2aGzW4z
nZMIXa4FysSrMJH6Y9O1gkyDdFzEg65LwCkm0FAHQFuY5/J1/sZvDj+Q/o/lotZNibhBhTR0asfc
s2EpzNdm8jIBNALa7VLPPMZcm89aswMFEes+JxpIzZrWKWPy+sWcupqh+Aoq4F3dNVXsSCG4Yl33
gO31pvyW0xRKCEBozXEQ/wIFcqp9VPYZ2O+UFgIVYtn885F5BPVzwtN8TW+AmpzVMKVFPoHGU92y
cKemIXOT2LnX2cSmvrnsBFjuaW2/RBx3iquSzMnb9cW4JXsts2zWq2uBVWMV9q6NXJuXbTRwrxsh
NIlsZQcnQLe2ooXiDXIgnnn9Vc3mvzNAuLYrRk7e7MBnZglSbOhG8r8X2LTlOAI17SPQdbyx87vs
fDep4PLFXTNh654/p9Et4u+uH8zjfqUHxq+YoEmwD5y8RGBiQyrGiVW/muBF8kFRNFxgUkBFOLYb
C/drauwgWnIfxDpFbqT0tPr5Ord4EhheeGWIMX0weK+qzwhuixHa/P6to84eq5CLudgzsX7UWnHz
lb3PKp7l5eJGVlRNg8hprRYC7lUhuPIAvqLqmBKa+B5uN4oLteqlzF5eqXVPSsO2yJ11FTJl6Vli
WL8QE7kSh+mfcluw8FVRFIYZ//iU5/y8lFw4xr/8jyLDwwMa1cqqlqBx3OCAHpVHYJ+rDccfGr88
hyhCnlxsQKJnOn5ohG82h2S8WYPtmZpwvTfmUeKl9Bc8ky545LM4JuiwOYczfpGYK9caH4QNitpi
2+mj6ox8nVUVWIye26bWGoYy9RMpqkvhHzOhV/nNDeA82QbWzWRicKRUQgxZ/oDfI0HNLHXPOHQ7
IpoW4WPS6NuxAmLE3QgirZ0RGNZVlJHNwyag8F9fChwhQlHFs5JnC9bVis87oKkz+OKeN+k63KlB
Ggz9NXgU5RkRLJHSs7gcpP+buArQ65rkSBuP/PL1GSv1Ia7+D3pMb2u/i+e1ML9AfUS82mc9Z9TX
q9CLp/0gL57AtlSJQbWhuU2tDKr7oknXOaC6W0gG6c8BWnyh4NVjhzvKynu+wtSuSv+gmp6tPL9O
cW2zEwtAvuvqABG/rJWwCZCt+H8zrVIsLNLy60T+y72GJTdw5aCIfskH3ID6HEg2PPIOsrfai+Wy
Usc+jta9LOKNvMh6yEg/g+6dB7484k/hzvIrcSCWgTnxqJlfwYv0KvnWbQ4tI+6fGg6DRXzl5CHR
NDPRbSvl540AI0a/PGbzkrFdGmeEjJvo/ymiHBBGgdf3PirY14/Y4PEY3ksb3JYFoH5CmpAZm5i/
sllXH40J3y8rpz+ECEIyYT7fSFZfC+8LMSkaS32AycnSQr0343yqgvk8NuNYdEs0vm3gLNzdiNP6
3ffuHkrEFFgqmvXAHa9wS2F0VZeB6xJx6tgpTH9nhnGEZ3oSNFZJ4milpjTWzXbvxQP/3wb4R0Hz
3mdnUlFeneHLkWG4FGgwT9YOeC9tvaT4HtUuxbWgHfqMQVpeMqSzAwDM5AWUyyDcb5+KAnvHtuvQ
4CmjphKY1I6gyIvU6EdU3ZlWtSYIfN6X09W1sBxsoAr0mnV0Va8xhPs4DNzH/6JiteAqX2bB+1OX
hrDSlm+MnFkdDajn37V0yvmBUXgGgnxrZGUGk74tT+tEh254tECN0wl/dnUQ550rJmWl7lxgiOiX
aJvAEUKSauHi0BriQXu3HWk2QIfXLqCvOiSeQypk0bvKEo64l2d76o4yAjGKuT5Cyizeo6AoOJjC
wg2gNYRzpY+TR4ZgbvZdzyH1dLuPyG1WK3SSWJa7sW8OKD7ALnbL59hhBZCNWCXuVLw+mpcLAtyv
+j4gvEVGbD0fZ8oAHNWWizzeqBlZTzyES5QX0GRTd5AnwT8vuWU5PBbK8TmVhwyLAN3XJyfZvAvB
T6tUe1+LFfOPQuzncRnuIo5DuB8xkrC3W+P1K+tJ9dvyWxBdQ89wkFIcvXfiK0ivaHwFPbnLq/mo
xHegQ8KUEj6m1UC+41gUhK2x6g/HZYc0UZapBdtcd6FQVR041454uUpqfG4zZKTpTuVj9LCJGaO0
QcQWd0LqJM9tGC6OYf0MHOPDTkJHlaVrUunCxFPFHbqfnewQ2MusFpU39zcJKEbigxs+Xyafe7N6
16GroQAyNDK3TckAzmnNH5lDIZi7umhztyikvJ3+D8fC2Bhu3h+c3Y0ioiHx7aDJLgdbWNpLerc+
XLMDwQ4ArZqylun7dYPZWTQluoiNTTHa4am0ep7UZjFbHVQFRjxylr+NGUKPSVobOFacV+gDd8oa
PYRWvKLi0knhrtOPo0EWcQY38IMqSSsZzTxUT3w+C2zmNlmC4CfALCK7XnYEncIVpbJSCLnkYqxn
k3ONw67z6GH9S/vY3mXc7sfrD1y0VMJih/S5HPV0f+79fvaKkNVxsdWaG6hd1076NayW/wOKVv96
3lHlJSPb4S7IO+B0V0QLhHG//Mvrwr74WmIU1TVoi37fq9LqSN0h3zzWmmJGgSGJ76N9IdbMA3m+
1Rmx+Mfw3HKFS++9cGUDS4aIqeea/VgMlCOrMCJn4QMY61tXdWtw0QSIt+bvKosf9JtvcPMCifBD
uft9PlSd9fENRD3v7JA/fgow1YI0rZ8D52lE69/hTK4zy0ddIgalAnhRkwwM2ae4iMBCdjHwRbVP
myRFFHan0XmksKhBMXgNoKDJrXu1wJV7R86QLcVOqzIJc7Ros5YxgDPmkq0pSv5jihVT4Gh/3DhC
RHlGfDFWWg56Ye/tylLxco4sIDjXX54wSApcalbAtao/mODBR7EmaD88gs6fiFbTYXiDAOgoxbvp
Nrate9UbQ3j0mwzOP1hZaIh6wyR9Mf7KyCoQYhr1t7zF5tykRqF7h/XBS4tlUKsn0B68kAvTtpKr
ImY3NB5lxasF5moC+rKCrFq+tVLE/d7iR9wcpIbbHVf2rfjW3eLXObReyk7ggqoCR711DtfeN2QM
cEtpsg8gneE3p7fdja/3pujS43t4w73SnUgnjhUxjcNuV2Ak+2HtJ/G4m++naNE9Maj9ymQ6o0iW
cyEG9pza3SR/bnoJ65nk4mavfdRhqVUZkDP2oVc3IoPALvmPw6o2SKxIovMsuZcRkXYQIHMyjhqP
GRg2TVvXnxgtzK7uOlFZ+DctEv9L6iJpBqJhTglbbcHOFXpMrytKtXC4bBtZtaunO5U1GuhVyRB0
1zvUoc65MMdFeQs8//vMWVzbQjzPlQxcaj+dKH9acyuPaAePJvt6Ek7rjpoJbcpeekXANoAHELO6
boRGWCe5aQyhOHyK/FTDJ7/b9FobIju+OmNHnIlg87a2s6Ct4s6doOY6yu0GprrwZYTWNM+N/uE4
OTrAAumOpHG8Mz1z0EN3KnNYHzgn566CURVQkHWvTFrVcnVBgIpn5IFBxyDTePGk+VOfywRWBnGo
NgmQbUqrfx7b1+Ri6Kp0uHKLoew6Tgnm30VOuzfycvgaTTQ2hKhu5YqXaWBaqdd64+6frY/UFsHj
YXw8ou4EFYu6lJYHZC1gcswIz/66jN7Aqpin+RDSOnYSRUcHXJ0qGzaltt7K2MOMC2UeyiNTzBLV
8qkxD75HSM+vHeKBSVIFGrCElNHub2mxks+GnmTSlxSsOJ3G/XxdhfsdnWn6rWbyoMk+T3hhHhx/
WjShbRLAX82sQS6zfeMQqAlvDeNfKOMYQ+qSuNPVjWlCRuf4PQTYWaj9oC4gHhHdnPV3ndd2mcZ9
D+/TCUSR1tVJqkG9NfdXvYeN9F3OOHLm4gSLSsqg1UwhqI0AZ9/2KolGmvKbhFDuo7eK9DTPTq6T
59lGxX25pvVZzx8PysQH1xBRnmhytjrAypj5BECE4DZhQ7PeRCAKNk+4y4zfKuKAwH7YyogDVl3o
TlWH/rZv2WtEyJYAKptfGCMukj6Z3eELJOPxoSAWlf666nh9aEQEB3Z/HXp8Ahnafa8n5+oN9stk
qC10FUDp4pMoOS+n1wF7nr05YbD8YgMcmNsjahmhetxUJjAUC7EpZgLa/Fl+lVXMRtbaONf04dFt
x4Lpwpty55woPeXMG8EcuffSNmpk7GFhBVQsrF8QkDGmsYteRLjeoOJYnuu+RJMNdYs6zoBawumO
FYeNi/psRL1yCvAtNZYS4OvWymYrEO6nOa/U56QYVUGVbXyYj+CS8Nu8zj/HZdiQ4/r0hxXQc+HM
LaiioUcVDsBnwR2fZhvmCE6wstNddty8/IGOXKxFu0FbKZp2KYfVagNTCq/oae4o+2zfGuaoHaIR
2q/XR7HI9qRnqFS5D4atTneBVXyObPFZrTRt7rZvjyD9TItdFxrG47Mwwd9DoqTjPRODCpFC/on1
PNkkjbDCzcPaMPUJ3SzwjtJeRY2WDM7OzEDMXuoGJMDCSjgk8GuNbI9faFa/+ESP4eBfenJ0dw5B
iO7PTNZiMgCGhFgDhCb2EWt3apAQWZTrhmA4llbcDSTGYuFlluiDoJxov5K3hf8AL9axH1swXwxb
X02pNGrBJgALOFqKee0wsB8nQaj4qRgCK4p3LhxAop5DtDuVyGCUpDgWIyPzHsk5CBD0FyIvNJFv
2DnZc6RgzF+xU2GXoc6MTTO+ftsUENb6c76T5JB2vMsZ30lIUCTCNa1KCrAU9HxKV9bNpNuKSpO9
2QtEOZUD6iTu8E8laH/Duer+s4cIEw4yOHP5wC46WxbTbW4EeYjA15J9bV2UUFfP3D8XAIC50gNY
jPfCdF1libxgkybwo3YT9CCI4Q6FwCGJsBAXOiY5wWK2j15X09xH71oZbZIQ/pBRFFBakXNUfNcm
lWqJToHifOtXiusUiHb6+QSF6soe3D4Z2XKP4JVixwwg9iJY45KfrSRuHgpriujSd5qNFdJ++hSu
nqNZPH+Qz7iARmvhdDkmX5faMJhuUoMCxM4payuI1QbvFZqtLwP432b/uGmsPK/QQYyOR2M4ab3v
dIXoHbIKgBxKJvThmaQv4RAtv2YloisHazsQ8F1vUmycAGxCEDYjHZfLpNcjDRQ1DRD+T19KIQba
r6HhP/DhA+sjzoZB4yrhYFle1pGTFd7nNK/53Ik+/4A01j+NtLlhv84GWyEFNM8uIizR0xBwAq6n
f5WeVhHT9tS16cq8JxnOnmla9YZwl7hZy4Pe5h9Mt/efNHyKp+NsB6IHdW5/QFufNuJe8kztxmL0
qf/72KOAwYXjuxneogGkFw9CpmLjE/wwdhT4kFsWNasK8q1Q13RPsGG1DZyH04aNfXHpp46zBnIA
oNhgA5GZTRUoN5XVJ4diSOu4d1s1BeM8yT+g1Hvo0n6I5LCVBLOAPhP22/bzPRUKy6EucreI+ME1
ewRwzlUoNEhV3caP2f5bXgzp0fXgaKQ/1xVG5BAtVPo6KhxCqJDJ9mZb/QgdTQH8QhvNjXOc8WZP
6xTXxobtLtlpwi3NP4C2aIQgW+4Da7zwfrQd/F6+CDa2cpH06tm0hndb+hztXYNCgDt6R47sTq6I
pVKesLTfcDSaZB0OJJQK43eSZgRIiUgc+R82LLTaSI8HXQb2vrK2B9yRycoZ/QBfBVNujPQUSm/i
ArF3C5t0FycOFbOqieTGu7TCnagIn185FogVR6Nc+RTev2sYpMFPJSzoUcOk7nUD3HIt2jonHdzM
BvZHSlna7i+dPKQL+Oqrhfj+ce8Z8lsreglivimOV/Q3y2JWq0UZQ2SCu8XFe6fz+XzG8Z08EQbm
UV9Ra7+KM0SGv+wc9Z/lzGZaUFW9OPa+Fdgu587kTdky/WTT1PtgP9qRe4hFmIvtP7zFWbqvCSXa
U8iUqO9le5KWM7Z8H31tIvKVhxPetUhG8D3lXzbOmg2MN16Nw1OTqr4RTOD1EwZzhvrGk8JXxAkG
KJh8E8hiiNWti8IYKfTLZ3inK4v3+Y0wb0dI1Rk7cHBox2BxrA5eBIB6Tj4sdXOUnlj1LdTYKcZ9
t1FeV1QSZB1mcQgVAx57SVapgST2YvlNtyO5nh4LkW1w2ya9SKiOozIhl3ST5jHX1WEindBC0Dqc
6CplNb5uy3pwGNAA+IX+6UM7prpWlaiopCEy3eeaQzeDtmbCQyvwywAzpEY60HMdlAhhevTMJkht
aFY8UX3WW6gKIhhfgGVpU1xzA1N18wXu8t8S6fh6MOMmj3rQTWnNwQ1HIhFdmKbPNI+C2HWxXzlH
qa/PW/D/JeWw080LBZYBuw/cOXB0m3Ao+94GsEbXzw9INS8q+7DaeykXBI8Q8NsAfP5tNH6nq40K
Hxe4KGbNjGcHu/hPKvALa9T7DOAlXRQziFkSdBfpnB/UhekFnpMLwZU8yjO4/SwuiJpe60bVY5sC
bW2o9E9HSlxzZFgahY1mhrG2lBWRfT1G0WAMXAL4ySJWyNonw2a7FLJ+KN4yE5nku2vJjoOUKjU+
McPW+L/RyDudUPFxt46A9f48aNsRH75KkB9M1gUfA4I7E+7xQKXee9wcExFbvag21YgTvVMn5V//
j3SDnn/q+6PjaT7OoIx4fPr9SQlX3jKpw3ZvgxOPLUrKHyrEuytTjyTGCrWmnRdeFK2i/MFhOgft
e0GHu4jvY0gt1k5pIOGIQHYQjxAzyBlWKL5rU+fac6LWUVNs1+gz8ucDd34lXSPBaJ6UqXUAT76z
f20tK7gj0sEgPvQKbHVaXdLPH8It63jfCdibzUmjfBMTOxzOTRrUL/iLjq7ulv0dzBiNEr8YTGBE
pTMvMXicDoziJOAUgM5xpYIzSWzGo59vLvuTUVyRl/e1rh8JljqWADmSfImj8pJDUdqjgXzSYLrH
fEBm+l04aiM+ouKz/EQTXGroEMts5TKNnV0Zfl8ZgM4wcVvloDk7YvvRKxJQTc4hZdRDWbd3bQbS
Bpi6iG11W30q+CfOqGr9XIzHKnlYZClfqiU7Kg2TbZipvcm5Gu1NPKPbcW6tkrK5KdmnUbekQBBA
e5d2Y6GiPBVeS2NVbKoiBgqHaSmyVB429el1+V0VMRe3GBA89QEunvAr+qxYfbXKHqAKYKAM/kHF
e3e9DjVJovR7TOpvHxyyMUzxrmvmjuKIlcLbN7NHve63IqX9IYZEWmoAVnxPulYEXCgSzv7o2wex
ti5GrO5IUqK0CSL1ie9YE//wnBmCl85BVcAPAkc/JKCAZU2MoUV+WtVKLvZhnPbFC9AOP1e0n7JH
9O6HS/b+kE65uLGa9pQqYPEYIuPp4WJycQRKwvR2hRAS0GoCZVcug5+jtcxfj4OjEzjyaBf32ZRG
zvpnaj7ewnD3k0WtXDBqc8iEsrV/4I1GqxxdBstwgO96/vx85CKBtgk3bhdOj+4oeVixS9iqlq7R
W4o6ku0N0SqS2/YlDKooA4ya7K22W0LiKpJtz53oaC8aEDBSWgIKdPv8a0yryNpH9jY7F2AadQiQ
IM/Li4PLVv/8vub63PqRdZIwDhMuacc9R0i93ieJjUwEUFqwkTEqVidc7l3wgMHHjWHr46yfLLPE
7ON5kS+B1SfYsk/WNU1yT4Gz7l6WEYBJk4keXDMbtxnBRfSY0v5vyz46sxn1uh2L5HuTpAbnve0u
g5/1bm6vWOhTfPO4YxrhEAkr5YFcYPQyRD8msIrnFFhS6BSgb1qwwalxp4CTg3fWoAm4eFxgRoBz
t5xP+FeUnQu5lrB358FihHbpU/4rsazc2t1R0QgZkaA4c+Mt+DYXdLWOYE4PhThJEmAsxbJQfKbQ
Dreh7syM5wUC1Zidp4iXmHXpAG9DtGmiNCIuyMUwQupoJ5kdaV7a2m8+pUKOqB8y6gDz9iJs2emX
fw4CYE+fpBhCJN/irM42gmp7e0iKCIuiuc1K3V7uO/USX7N6GJd8ik1czhxCYzh/ol0avme3rgre
f+Uge5UqpHcnO5gSj0PIuUAjwMXE94FSHxVum7XE5rwBXoXcdsFyc1h7Qz09k+n1w8opSasim89W
luQtkEqIObH9+9vuU/zvhYLmCSIbu3wfqHeFzyU6fkjt7hm1b6xlGp997oUsw7DPOEu83Fub6Pwk
URaI/oQ2JPzwraqQ3tGDRNVP+fMQCU4bIGeOcxxv9TKMMExjOI2k8B/rLGCsb7or/2rf/xDgR3Zy
dSP/AY6zuYokVhUiGeDq4V2WpZWGOgDBOAZXRQGfionUHFhWUHFNAMU4hCC3yYoTvxRhfWz8vZjy
Cppwjc+KJdemXz4gz6GlawR8vYN2TV+VQTe2i0ImfF+33nljzJYk8CbSDYE6mn/rj65rUljzmZgg
wwgxNLetapJPxS5ogreNRVMx+pCfZMvhCdgqLzKSU4s+u4bKwsPBzklgNPy1V2VesGdQXNqQsviX
L9aIOlcKsyJz3/hyAuGNZwIByXQ+B3/ZAbZQlISAjywF4z1zqrrQcwaJiGFaSLKqKTUQgi4apbnd
Y9kjVoNm6XtupnOlvF/2FxZ7R+Rp4FGLQBhvf5061nxwCLgar7MwpvX8Ad4WKIZHz3YgdVD8JMc2
hnw1+Wke+8tsZimw2IEl9E2/usykLiEa1H6SSqqNPIZqGz+Ch/0z6GmncLiAstLBjDz06Rmfd+o1
4k50AqlpIIdQ61JnAV311UHHeOfmPUam5S9PrP9jrq5U57b145Vt28pZUNMAiolc0kMasxThCPGd
XZRVcOWeUJRYi4iRPUk6FdnHXJWYFrRVv7NODO4ELN771rjSP+prHSPCJok5altVeeedyGRavpA4
3VBImf1Ly6myPWNb8NxlCqlkUxN6EfuI40NU6L/NZHlnyxGp590Gf7LNAJMcknnV/WGgdwBfWebN
FdYxlCqtwZaNf9O2RM+5A8gusDGCSQgWhyxsO5h+qMO1h81OEaHeV5+tLZNBudYR4OV2M8yM/Ufp
jPY0P5WVbyy5AWAGrsHlqsSWWHvntZ513SQt2+DGPnEVbl4qvS27uvqkXf5/Sf7sigGOyd75HNWr
6slY0jDzzCFJ22uQ6LiPB3vppLBmIwsawMApogNUOnfG0D0fcPYaTVSsFOfvW+SVzvpXlUpe3pWE
D739DpnKCRO02gPEu/7ShT3IshMOImkJm31+jc6zj5Yr6dXkbGE0SWzAMhs3nTIROtrE9t1++QnO
C1dYURQPr02AvqkRO3p36JRspxwSDz/02la/aqz1TVkRg0DG3rONf/wCTkwEDIvsY7GRE9RZprfE
vtvSJzizbBvzO0phxwIkhVIgWFEOAByZwHncgnCLZq2yHPxFhvg8jGw6TEEVOILv12obGelD+tdp
MR71y+VgkkgdNEB3hBhf4bs6YVygTSbK0RgbEPu+zgLES7s212B71p0loyAe54Zska777+10KE+o
HbO5jt4IB1gNwgycNQ93/Ydu0z41P5qGVRCCPJlil+MZrsYyePe1uXWVgjurDEkh0oJx1PSp32FA
uQwxgxQT4vC29LZUjmDgZPBC1xhcqbuoGVDKeWqJuJXnXAJHXW2kEWi00bwPMxeKUSlHRn3gRzGM
MogcskUgn6NLmAN0OV6POh90KVRslxbLU4OuIDC60qxT5bt8LrKKPVpbYQ+kxQce1M5eg+xCotoX
MVgveM2KkAYZnCEwmlZz4FfHH7/GxjTjnWWMvgDWYzBuMn09b0ycYQ1diOmmj6jt0E8u56LxcuAr
rGP9WzZOzHN4zoGg8HqvyAT0qK6k1P4tdvkMuNcQHyEVES150SVNWimQnQPLG27gU15KEdR0pxVf
ZRrIqCiQvFEDlAuwctISvfslsW9u7GfLW21i8FPui2GjI91YWSVDrEcrSyZlOdubZLAuKGrKbaxg
gibnRVlyCieAQCpmcA3YiAZdP4YJ530L9wTiqIYQDklzzy60qtmU0je3L+oX4/Y4TU4gpCOm79I+
06yj40QLwqSA8nq9TWIfXjOIBLJ1W1/vtO4SeAtb/unvARfpMXQKp5Rcbcjq2rql79HpjoLvvWJr
FCpC4bwzKDT9RjBfKSpP5cz5LLvNZa7ndav/APz+mxaOOH+3xTJm0MibzjubJdIwLYZW2YfUgO1o
oRBM6WIAuGihwrb/s6hw3duBVa1XPneYtMqzmiKpxjhHGncxnJLr5h/cUqPNTEXgGBuDPYFXWUJs
H9tozTaOYLDq3yaQ8LjflZwnqMYpA54DzzjAAs3xWn4vrO1ZPNNQ5IVPmChDfWVHlKhNMj9TULQh
D6jFF/anE7waJYJEdx/NvcAbtHpu0ywOV4Uy0R8ZreoQebGbpA7T5zM2Z4qgsyJrt0m6/QNRASMj
yjMKbglvY0UQdtrWnMvRa+coVRm8b32jlW0HZYAo2Kly9Oe59zBe0xF/REqLiBPoVoMmm6je5QFd
6inxH5+NfVTnhe8BGb8zblbGefpuA8PSy5Nu/s7qtJG5DhcSboktj9a1NW53tkP1lGh814NfiGaB
xImKz4HlRCUS0+G1+rRy4AMTSSbNWII4YaoOzSZKHtg1xzdyA3I5l5gLf2UqZ5Drs02NJJEMr1L6
2W8+JyEFr9UQ2RO/DbHpVGi3Qy7hi9RYQpXKQDmOJBTYNkmZ/gdvnbW2sUQqoWltboL1ld9POM9S
+qUMn7nHTRd3kISHNENnK83AJmhJuhRfWGh40EbLrIfKEkY35F+RKZpJ81wV+UpQt6qJKmssHWkj
hymXndTDSqZk9jfvJpga6MMkk3NHOS0Oc+WGO3xgAt2ZDzE4XTz9SQgcI5Z2RdCfoeNkRT7Ujy3j
qCXQP6z67EVltH/wZO/VOZzBpqEXONET3rjoXdSJiOvLsZ9Ikjc2tIflI3ks2dG9mD26InoV2TsB
woNlmJFNB/MUQfOwKIGyq0CoTZ2iJ5XxXuhvOmHqces5chGpjxHVqDj6c2vfdIeWB2nxajNicTVm
J4ZyTFqdOPZYs4qaHFHiHOnwd6CxVOCs/Gb1e0B94u1huIDM/2EJJdnT6T+aPG5IOCPg49VmGC8L
MB3MjG8/rfdSGn0nsjBKASue26AIpLnr8zQlPMc4nxPmIPZmN8L+DFogqxszdgPB85PoBb1DJFz/
fNZj1V+aOU2ADczuri505x/kB0HSnA5mWdAkdssy6mjNK2NEAPMHInMC8JwybDbhWPp+/7E4otat
/RACm5L054/hBP3vMbObB2JjN6gN8xoLKaf/tmgyUjbBzBNgQGCzyuVD0veWkaJjPqO5rU94IzmW
hAydp5gR+LFJQ02DFWx7oOEcyY05f/8rCAh3VeofBtdPMzFd2cnjGk3TvuUwNqFimvieU7UGAQYA
LEzQ2PyCvtEaUchH0NGEXO5JWsRcLrNU8N1wy35jMYyb1pekqgXdWVh4m0Gtik6851al56j1J8VI
l4xF4Ond16qr7v0qAv6RyHU+n324jpmq1n7PmXYMIzMPDrrJgG3sz3GO73H7eKhg5kBsMK/1SlVP
4L2du4kEA72Ukq+RIYmdUnkLLWLgYFonWOPRcfkO7dSzFeqXeoSdbBaPpYxLPwg/zaobjIZaA5xT
YM9ru/jXxAvSaSyzhuHIA8U/2tui8KNIGW9BRs5F+gZ4zv2qXcVvIRHKs3NuIl+KyjaLmFm9WuwE
zxyQLM6plOLKYabQ8w/pI28I4MECHFmWfZ/NftdyKUoh7IMp9AFkX4hBqrWqwApTbf251qL/3673
Cz96i4hPW86s0RK0bZdOaed4i/757/fz3DziHJG99f6LGqjdGxcmJbtzZ38alDtDG6DnAMILhEdJ
1DLkBgn30KfK/1bynErys5FPoNgdEB9JWC8AhFkhg8APovVeHVYaOlo62CF9uVLwOf53SgVcXMNc
Vuh3QxN/gyVBa8fAWuaL1PP7CFvmX+e7C8iOFp8bmu3lHDM0ZC9GA6JYCvab651nermSVbDziWc4
T594EaCqm3w+4tvX6h+WH6GYRSNg5lPcIiQMotXuE8RS7VMLUi3c64Z6M0uvNrjxD7MDOKa0TEFy
t8ohi/h48YuRvYNDx6CxpQd84D+0nQqOuxvyE8Mo1I7N9L/qRojOwMw/Tb9wCC6VzkwXQ0VrAjgQ
qurnjf7FL4vBXlmx9KlhmTqm5xD8L62DOeVmP6pGwAxGD/Yq3kWn5xlleO6tX04HlH/9M1NKHaPC
l8VupOblQeFlYzLJMFsFuH4eCRTCbaFvf6LMLBNVVVoJNJgRB2E4BTqeE37Lvl+Vrw3ANHzNW4fu
ms+39eKePoU3aJwbHr99h6eZb2Nfv8cfxdzu0FUopoCWsO6lbajPcGw/hlVhLwscDGAN0v8BseW9
5LxW9hFiXVRG1zEucSV6CSjTqrFPOZwt9St1QG35+jU9mpRbJPi98vMZgWm8pr8AKsdDR/1I1fvf
+L/gv68GYzuhIFmG0gw+7+QOVflw38kC9/O/8/lxB6f1qK3wsk/4iIOuVN5eTs3dw/Z+EMGm3ozO
yKd4+DTq8qq2KEwF+giDo/MyBYs1ZP9wkxeWKdwJWp3y5eaVMUJtuosuUcLT6PtsnXfU8tkJeanK
+xwbyK+ZkCILMKzgsfhg6jB+fd7fvJfcevVmZdq43MjcM5OnLGNXkNERpKYTCqfSpMhNbyLAWtPf
bu+gntToFD1s4EjLsK7SUlHFCXgx0Gx2Vdhr7ikFsKN0quNoKrVzjU4eq4KEOSFAs9T4GoH2cuQV
55GJgGF4zQs2JYcXLuaQxqtmRDVug5VLt8xYZn0laN3krZ/EjYhiWTpYlCvnwWsJ/l3fBiEKY1IS
2rSbMBjTANZjaQgUSFckFBW2H2kSi1nzzpcd8o0VegxLgSGPDtBC906y9WDVbhb06+SjrP5MfRYc
xvW8V/QSuA/VdFVllQ4XY30Cv0gdJFr3DQpe2rSANZ314jjhMbp6AYVaWdabdhUzLGk+Ui14mD3B
hmiDkxTB5UTTWWbi+ETG27w9bSUksGViyUuD7XEpqJcVMo4f4cp2jB7dggnW++qYFqsmF3EA4p0P
fFssEWIfcZ3QxUxdut4mDzZhC2eeIqli3ZOLswglKV94TciFfefgmHVnUG455Sx0yMGqpduyBuud
JNaYm0Ys2bt6dG4xezsan/xNF5CgTAjcPUov9TxqsmE2eNX+ZK/jiRpVLirtJUoTXWp27KN5A/JX
hJjcfCqP1nIkuzjSrK6e+ZvsXsYYR96X+5zdq9VcSMzhCFReHWE8UgBqmsdM6m2sxWU1tAou/nIC
H+ajbgcEFbKQg2WU/6sy99G2zwdTnorTdic+irYLKquhK87HZEDWvXIVZGYfnkmVReFVL7HIH792
yztRIkf/WIjLOk4xy74bmwksoFZJrC4bv1zm9+tssHbilrc4N4Vbus4mncr2EmPiaMDVTGkpXvQO
M3J8wjO8+cCASxENrc1Moex2Wwt/erwVk61/UYA+TGdx7wUQsp25d94qwpLHAjqyxw/MISAFTuPv
ThYkyHxde3DrHsQJofrtqsIUNtAC4KjVnnNXMQu3FmzZYaQl+hkzei9olvuDDxjpGQTTDw/U+saa
ub0fEZ1vaPMEX280rqb6v88tKHB9t7BNm0TkktgS0j0CrGPszPM99k4yCw3+SwYXYy6CEDpoVHpW
NoDI0DQ8zjusPGTvwPYVoZDWYeQ77fnwubsAqn5aD+QsPtBQhpH3+ra09jMM+M/RNVIah8++LoVD
A6XkdV7EdkmdWLhyJUcMCPB9tQIPjuA3Ef/qWENiNou98C+9oHLti2zuLFDVl9PQDmxloy+PoqKh
qFXF1j7dZOzRjj9txMNw5byS0yDYz8PdSey/oBQfuyRa36d4Bga9Ry1tMH5uba5l/+npxyQWxVSf
Ug252OeBXH6VkAha23GCkQcJS2qf9R39g0SDv9Yd8eEp4FDSMJDUXu31bpR7NTeLHpJdKU790N0C
dhCNIaQ3qoYDRbMPLiArROAcHmwGIPR3BiIJj+TbxVJ38O+P0/IUApy5wdWZFzhBgwkp5UBuN6/D
uj7JMZiIAHR1T7ro28mJOqFAzzzxXY+l6r2i4i6ez3lEWL3/Dq/bLxBOX7FJk48ibgJ1Rmn9Ycv9
f89hFYATctX9ixUlsls3EGSoYbjQ2FkULgSvVsaVv5xZhMYeiVvjpwnDGpMxkGJvJW9chTMtn0w9
q41ahZ5vEVYwNS+Hb9+q6Id6UK/89SVOXSzqjq+kUoiriB2BQG85QQW+od63oByR3ErH2ubMXYIt
K7JNl05sWtZis+jHJo0BSYKEeM1PhIEAUTXuc6AE/sLIhQb8bQNv+TAuB1MudMxk7oK58D4ZX85B
JsuSeD7JSgeKlXwAFSTmivItqTZbxfOoWBrmBP/t+xF4vWYxJ7FK2EDJg7vd3b8wmQurtp38roEI
ecCyqb927H/v//6LVQKzK/1v3oCkTVNi4k0z5PBkdQgGMPKMYwMuifoOYK+y846Wghh+dz4fZm9M
hvEyX3r8ZyfWIR2LCyIctrm8JICOjofT6D8/XQLlJg7uVklppDbbYYmH9G37Xdv//KoF75c8Z2cc
3SgZFawncy+AvAxNSpII5prq2QFD4WL0iMUSVJj74QtKvNRP1jAKcOzbfF7hwqRlYIFbNAYXp7ZK
PeA2KtCioIQlxWfMDoOpPgSgfz0YS3Qfim9/piwIogWRVXm8ZZXFc4nz0kfdPdJs1KRd5VUzGXdC
XhLulOLxh0TKKoaRcaIKBPPEgPlPocLKOHW5sIkiLiCltmK901VbY0Z8pgIGSTNt4zTCjNVXMNtH
BnBasOrFXz6gfLYtQaEmYk+YRvRa31KU4hEHoxO+8UjHmThy9nnZUAaynaTX7+WOig0VlDM48kvl
VtPOPiTnDVegR18Bc+IfKm+3IHCR2kE6ekMIwW52ca+CaQ3qUm6TmD+I1oKeE0QCr75ygbVIdCXS
BIgtiqEOQwaz+Wx0ckrGUzPgi78YCYzOBIN4oVpO5pcJtm1uu3yTLxK49Ebvng+nwypeaMdNiQpZ
jmhlIDzwkTrZQYSrTV3w+W1PPzr4/DYD8BGr0NESqUDJs5TxwoQrfzd4izuhC5tw9yRPP04pGdOn
kVHuP5g7seFEjp9m72ELYAzYA/OcW4HqrvOlNJ/mQxPrayqnf7eNQCOUTY1fZxi0yfcV00Cxhv8o
M0YNwygk4mAoEOjAT5S38rv1Q7HFCIH4wOS3++hstoaeiObDKA+tS2a6Vu5QEaZLRd4YfgG7kLZK
GdwYLdMBx9cYCAgulRU6CNyWkwoooN8PIo0+/j79nS10JPYPICxBW+5aPgp0YjODAipgGQcAVF2i
b9pmIJIvvpKqNfXPW+c5FodHODCmUsXV0OsvFZTfHWROW4l25Tbmjouh7Yuzt+cNHcy+bb7SjiSR
26+OWfoILBUdDTvePcLRqXoI/hJjms9Vrp2f7lbo9T/AI9X7j8fzK43HHufGEWDK3iMfyBsg7BFt
tYSVonLf9Z0IFk4Mk7fBCOVYht4TzLM/sH+r5cj5ZuO+2xpXKOhjBS4L1VdocC/j0CNvhe/cQaeX
n2ihUTdV2+Yg6HCNGjy6gEZHdssXdGskWhlpa4zMF21Y+YLmZcnw3OVNOlIwAnm5FksRMerviRuA
+6ybvr3BI6AFE7Arx6ilAeXDshN1PtdYwBKhCFBUyW15xNKg58kVTHXSzOmPi1tFJdK/qifbUyfF
ILWCOh+XvXQEvoPN1zCeDLvmwHucJ7Vj8BCs0frjy1GIxh8JoQPb/PVhi4Vm/QhRhPaipOTxA6tK
nSFC+TiZvzcCmHMlMTwl+9ssgzg/z6zn9Ym3ICATSHz9rR8esyoPJ/nNC66WkfrZ+mJClKJoZ6P+
NMIqR/1060J2lIEgT5UxkakkR2YGiAjsxPvNbuS4vLvsOVw4CJzZYU/1y7aW4jFYo0bCWVbtjgZC
0L6EZToLjajLOWzQF6lzmUOE6mer3QX7kx+SWKOHBrCR9To1hSDHZs08Aqg3BFmGnb0DIxNte84n
bcFuLFDtLQJoPYmrPs/mDmTmYpOcp4PlkEUV/VnGSxCAeO4WJiYcYnOl1q/+QGngAJwIRMPhozPl
dLDwgN3ryJnvZsCQvIEetuce7CP6lkY+rNeyDo4fJUKd2585jDcDOyYWhfhQKYbrkkvHf1555YLn
4IrS55HV2EdRljAXjadaCsxyazw6znRMMI6ZM/DfIyhBYqxyH82PYa/giYXDR6YoKc6iBHnIIBlY
/SfWv1Ez1sPGQCpzlGE26bUo4/KwGRXLfW4/hwYiSby7nIEaIpxqOOZvmFRrGGVGSSKBIohUFDrt
8DlFfBMmlcF1jz0i/4eJAAQTupLkv25ZQhJNJb7N/pNcne64apN+eaa1Oa+Yr1M0GfbuV40lTvkl
Btbyjs3ZvInUNEGgGoakhr42ACE2RX2B9PpD5AIb6Ox+3MjM/dqjwgoeGLG80Af8Sl9hOkPnyf9k
XzclUhUSEtpoSSKuoRyz0iff/y08vOUdokYBIvNkeBfmhd454xmR/JEwRXR+piKPjd2xwj/YcMHU
MvWR85HJt/HhUn28suxOYTIP/pogUoIdoKOuajLz9s9UMbpopJZaN09Me2nfTbss01fJUnCbw4uV
4/DY3fS1Q7Gf2BDE9OVDxLctEHwID0Mo83PaZsT+09xOFtt5B3jS1Mv8P9VHk43Jk/aAaxUMx68E
qLmIpTSDt6uhXasihjB6CzkHuXnB6u5SNHN0vFQdUwUyH7qgen2UuN2IlLMpHilP0eJmYwESMSqv
o3CBfsu6DvZbcvp0y2TuIhFVsOxVbA4jY/CZQvi0Kz0Ia5dQnZHEcz57FAaVtuIHKECrk41jsCub
lToG6T95n4Ofs6LtU1Usd4OFe27QSaMDEMBrjVLnn8g66h2jPKm9HzsqtGgdPQmntmhzcNdm7PCn
ZzvfB6Un0v4chsxcaUnuJ/+qbF4rbqhlshPHsSeGgb/x8yB8NSO/IHvSHwym2YGj26P+K/4FeaUD
eYmk5Cp6N7DCNFStjK6vkDoGSwcraeG9/S97oM7srU/osd6iomdZlgdd35y13orT87HcRNNDd6e1
qa0UAohbAh4xjq0Sdki09YfDos5nREoOTfpeiYVoYHrZ/COjBEjPKVnlAB4zBXd6cN1nybCakEzh
g5bKBkgor2FnwtcqMmw1dgqBd/r5SKgpCYzdTCKHYkfxnKIw92VBpjGxjGsdhmsVZ33nYy64FDqj
Vkm65VhCiV12MeirO1r3GwZXZqwgnAHe+f06OYZiFLiylbtIWCMqDm99PZKVT/Dkyt+2JR3UFObM
Vux62QSDBUrVQqQrwueam4iGWt6GeTDoyvpxkFLzUb8oTBgSoagBqLB9UyA2GJs0IjYhsEOBaJpB
8vUIoFDkAxAMHgZ9eSQ4Z8NcLiT8xj/mzWw4AyVkhHSn/RZzO8tNY4CIS5VJUcX3zSx8CSb+uqmS
O5ZCp7XmtYV5J7x0DOrx1iZU6R6xrUwjmUmIeBvE70fTzODBbgd9Nrrig9D4+bB9iokKbd34S4vA
CQXWkvDIhXH1qiutzvMTYGvS4PKoiacG2QstegTND/TKFdK0AJJeUMwzmLDk7mODBjSrEClIjtrE
VRBMTG/84KYuvdkGESNlOhZ3dhzLJHfwGt21C3KIGCngzscCfNLVCtOO3vbEvZta7YfCK42SWhnC
1olcOP3pefQDfjdzIq9vABFNj6J/eLZzWJnv1aTyXqBnC/BXeUBPqt0Rzvz+avyMFNXKjbEIX7aW
2/n6eykPmS/6Pg5Il2WhvhTS4HtUPKgKPX41L8fW8wRLW85ns5kTfHa8TP93sOq6XLA5qQGouhBi
PfC1/NdHJx8OO49IyqU2V4NbuWHjVibn2n3bQTTb6lGLRRmVk3I8TpjOFo8sJecQkZNgVkAT1tRP
fJwX3q/jl6noyn1ybPgEwh01dK8HG7lyX2qbIUwvnoKuyk89ZF0ubKZZfkjk/BXUr74wXd69nNRJ
du85nbP3MYXRd1h4S/JlszyeH4mmb6ubQgw2Eichr9V011+CUW7v3S+uN0KQD3xWR6yQ0IphGQX4
lWAvBs9PSfqtGg1l4ct1z/kwudN9ImUw8IgwgVj8Cvv5qK59hoqWFc5pIyIdCsnvSfJesEO6A7Mr
xQgi2Xo3tnB7vqST1fQx+6IV6FKkZsxLfsN+Kc+zYSg1mFoPAV1dDqlD6f0QHlBsFVtWS/x60uzN
/4Vzjk+95dccNzc0/LW672qS0Lv92wVcW0MmpIe9OiPYiNtZWD9XH6O5GeJuIS7aQK7EyH/OTxzU
ZhgxUc5x3jyy9t1vjIj2Rh1/bzudszqbaG85/F7kTYAgmunURLDPN56zm4/BUGq6BJEiP1SiZTIs
ljyj96kq+LfY3gMPtMQvwtgN74AXQhjAG8NSQBGbRvFfB3FbEKO2nTIOPR4pNgB9HC2gBL4J5+7S
0npOUrmqee5SalCbj0ObDP+H4CfZU8OnorW5N65QCyla8N2MXm/9ky4+vUaFI5qDas1nCBvRDnG8
Ei0OD3aV9ImKg7kSF0IrFx66Hkah90Pf9FtFVLMgYfMKiZ48xCBlo0WL/HWcDgUIg6jHzaK2SLbT
Rd75RYmiB22dneJZMO/kKG+TTVTty81KdUZCeFdSj2PfNH7CdDJ38bipL7Zh8AC0duqZsCxzKy1k
R4TrkwO+rOTGH8lfVEjJe4kV38TGOyiz9lYTgRDZ2QPIYqUQpnLhg+kG+/9mC+H3jsLLq92lZBE5
NmCMuDY3oAJzzmWM5a349HhfazK1+JsIOMHzxh3ZN2aduS4AKq65hkziaUb7d8ZXdCXtEq72+EhG
7h0Wrj6tDfjOvwn6T6/yZaWeGnAv4p6L9Rntz4kZlSmdfdN/VM1VdJHMaPGnGdmt4qBFIzTqV4VR
iF98wFq+w/l+UYUei2slCA7ExtWMopkIdohjr4LsdgxL61p0QiMOasMYGFWQN+jF3yXxwaxjEvVc
Xab4VLhh9h/4Hfg+7oXqTFFXYv9koGLplK3/fTSqosiJX5XTt6UUqs5nBNbsjBocZSTBo4Hy9dRs
/BfFKgEG/grPcGroLQqF3PZROW77oOD/5dFzjsOiKHQgXT8fm0u/6lIhuQ1v3YaKTkUFGENuP+Xz
gRSlGeHwBsfeHKGLljvdQXrIIxFIX8dcjDoXcznWrodMoedMvLnMPdGpVvKzGyFYTa2mROphAW7Y
BcTntHo8goSagEbWnx1OdDaH9eTFbR4z9PbDgaQin7rn7hv1y/3NIk5ySckaujcaGjsL9q299yEh
63SowXBExRBIXdJix3wOOWxghW7dtPkuJlvjO4ZMCmjDUKgyk5Es3TKf/umNGt+zSzmzIlkRYJ2z
Lzi24Noqt2qJgrWo8KmNcSMo/GuJBWztWjFZItFyyuik1BgCbab9vyfpf6I1WVPSGOUqS9I2Ynpn
q28c7K9D3BJsYPGF1HjG92E3FNMc87662ySaxwUrnKmFWHD2YHliK4rPuqOz4d6w3ABCbOvkvp6w
rMczyQHf1cZQ6g8QcJYhD6oI/yrTaVEuqHCK6lOxyykszAGZbJgC4X89Syj/CCECHEN+98mNeN/H
k2fPSzWvWwVD94Z8pUOqWpj5GOquK1o/iVBjMSb5EppohSDErSm5mqfBhNPtQcF/vXw/l5GxAe1I
mlNGpva71AVn1nDXS3jZSDraF6Mwc298WZc1lco4Xn6Kwdo8NiOPkNrdHz1yeee2VVnTO+QCLzI8
wGh5liL3q45ZfeNHExjwK3+NDH/sjDPpiAnBoGITmqx6y4y1RbnxXE/ex3jy9XuXexSlc+T+YIl5
toZFeyChs2WLKk39qbo6w6z02jK9aqGhyYRgYVu3aZa0yT1uqoYcS1F5Js8FfM35eg08nLu35uER
fmoBLyxRziYA7c/w1lhD0Oognv+wL91CRDDuBT/GNFbEzR0QwQk5DJzKPbiKqGj8pi47w4tNWD2n
Z21X9PkgHD2gOnEZAbvFRzH27aHIcmuZEm2tKN73R06MwHFpLlKjPAS6kuzVlI9LVWiF4EFrrFV8
2ilb6TtiGGQXjLZb1VUezS9LoGyDvGSppqg5nzaP+dgcBvFCZPUsCYR/6HzQ++sV44NNEZ5G/IqE
vVb4T8FI6nf8MDWAeiZNU9NgTXPqfB5J2YwqRtgLdvNQP7Z2LJKjUZt+r3lIFhgLTUMmswJNh23p
YM6UdY7Tc77/8TTn6iUY7v/3bwVLIxvtYAPnCS3L8RWs+RyR1x91ye/xwisqxM5BOdkzYacUK4Il
aTPxQr/ejNA/Z+HNFz7dVFgj4QjmT1dyrgYECWa613pOwVx0ZsR+FRo8v5znTbi0YgFDoOSOQkW/
jl+8yxZul3jpif23z134BQno1sy9Ty8ANUY+PprvC3AER8/4jKA5HY/qp/8LW8IHG0Mg07Ojfsns
gFRr/0//sN5HhsYBv9A/a8cq2xFxrHSv+YUxezpQkslxoNp9T7hgWm+cgPYBvpyc9w+vG14iywf9
eY6cnVX8aEyGAj9BrpIP+v72oOXRAeOUhHKW0mydAd+Vx6TFLyCBLcOW8zX4nEqKDjP/0fNig3v3
AaAXqAeDrLfXz+lbyO7yFGRMxXnUGOexvnYgzOeiqsCIRXsSVpm0HyZIlJJQ5vjlxCsebqgmnfI9
Go6cVbl4koSRhHjoaFaeSz6U5pW9JgJGd85DHf2AbEZkpb5fDk+PXCQG+SiTxNZ/td6qaKJbJU2q
uziRvuz7W9WmL4VTfYc7jYDRb4S9VWymxTFN+SMVF3flASfjo3qV+9GHkcR9wVkSpwyI6U9UWyyV
1EQ0TXfgDo/EZTeP5KQ6iVmXLGVb69gvSOskC9qlNxJWucNTQSRQb3LmxSd8FRWsvXociHBIJ4iA
ajGiG5UvUDoRXgiQ62yIxmrB9TjQ7CNagBV3xXZGkMdIGu/VlRG/PwqaewelgERpMYTSJpPO2McV
RocIT3GlOj8EIeW0SYDaJVMdlyB9KGUUcdqvtPfSPDOXokfclYLlNcNH0fXH8SUPwEamoyuq5Djr
g3+ndnrXV4COp1A3rDAnDzN04KxvsoXtHeN5j0gqHhSdB5QACsL2fGqe32EDRAScirnzbYtBEeFi
altfPyF3p++D1bZyDV/76EkiZ0/iFmllg+B1mV/zwiyR6ru6pqGbX+Hr52MiNQTkp6N4kwGKAnw+
Zu/yEcW8qWw2EbgceeaooSizvvgX0SWrb+JtkYvHHAstPBjQwhd/b89DSZTUarTcuXkxnvTVvNUy
8MRpZ64ZcFhxvSAyR/N1CqPfoq3GwEJjLqQLNja5X0vYCBwMAM6us0EYgm5AZ2X6JCAkFx2QTIHZ
eQ9mR3s5OCjvXmroxR9LbXvx5xp1zG8urvG2VUMMLi5OjYGj2Crj6OSBYv8TQBXocvdW0YVPq+ei
1C72XJOyZI946FCJkqOEUGeL7HQ/rTwfDOSW+bTdz43s8SorsT54PC0W8eIytVLeHKMNCPD+3lV0
rqq41DX+EHgismKgP0+OCr1rIm9xHWdvdFkIwDl9kSoeIFl/mAdZ07YIwlj7wD0BxF6MmeRo0tKe
loa5nWPghK2LpD5tVXdD2y40jRDisQwThddqsSMQVJeUrXuZj5wf6DifdOr4rHoKaTWSzMFAhZQx
9/kSNA6ursng3YC9JHdQKiBQ9OVUwonyyAls5mGQ1AD6QQez7IFriomkd1XxNkAgAj/h5hGy17rV
waF56OPwJXEdkWVpgfu+PTN5QKCpiHHSM0WqpQsM5NA78Hy/ASA07EwYEr8Pw5ZIr4wqIUHbOv/3
4kFXbmFjR2hFHNfbjP5f16CEyIrrLrAkFkLugsI+1BvVoILGNB5wDET03vO45AaauxaHOIAHcWsp
o8hnG8PCcmUV8XL0E52oYTqHxkZD0auyUx7Hk6sZVnU1ahXQxjuKi54YsdvYTHYjkt6pPkT0wVF3
lW2KrCtNklvjux76w51YWSSjT92Qj0EXNmrOgUw5rVEifd1z0SJyYjQ8uAeu+NqRTqhIyssSMw5I
pEj++7CpgeNl6tVh9FsyyuwD7MYrTfYp8f7mrdDp59o595wCMhn/lEmnPFNRSFyGoPigiXkCzyQJ
rdrOW589BQ2kDkN0Tjsx0G490b9e3RRuJcaFDYun2E/IQB/ftDZlak9oFQcBRiDS0JYwndG8EBBA
6r9rU0V8/TVRLngukruTK6gbyyW6VlOhBQoOI7hGY7Mzdcymfx6pbXWOfly7Cmq5KSDA+G9+QsJ5
FLmzQCmtwaflCMEXQKzGHFuAQs4INwry55nvZ+JohKl7LivPJKX+H7vLA8Lh3BTwQG9hPceAeAlo
Tdq3Fau3jwsf0wQ8kSh8eF3TrC18Q1RvK7UlDTB7dFXRLdUR4xGINvVqqyqLeb0XdFWK8i7iEcnF
gVxI+3plUPqr+mlDVHwzQe7Y0boZaXAqApKVaoWHt+tc8SWjbO3h5ccssA7jwK9w2fyLAOr+YsmF
058MX66e/gfKtxeqXBon+0g9k6H7CwZ8XVPIaRBrSPwPMGqDJM1qoovd53MiyQLhplrHw62YPgIT
dYVIoXRORkNqkQXX/Qp62oaXzfI0d63lge6mFDPthQZTz55EaeOKNT0lrCpshhZGDRyD7kmLhwsl
Lo8bBFtd9Frj9ADt2I/nXKJKXZXVQy7ozP9nEFhvqKAmbFrZLLBvVDQROgfRZpzK1sckwYsqR6c4
Yql0dM89Jgt4YZ1wEOA9+HQtu605TZVwdL34YLl2twjEjW7qeVY7/KDnJm8YGnC4S4/NI5hiFMQJ
kTtUGTgeARNPjsOC2pD37jicbCy3Z7cKgrch4n3Oxn3TBynuHpw5PMdHWCoTBqUsTRwhOw3qN3Gi
6dzI9d97CuP8LOf9RBpvDs+mX3sdG/H7D3D6GyVxS1Bj+qizlc39F5Ja2FwQRS+XJu7PFOkHaIgp
jwOpt+55bllQ9be83ogd0fgG8myuZIsVh8o9gnnX9+KmqVoyrBXG1jOOEuebFpWqok2wlJr8vi2D
jzMsEUrOe73rm6rSQrHNM/amj8afKkGGvNRQTrUEpmgN7EbqRhLH/CiRIQr6I3OVGYcHz/n/XWMW
xXgQSLtaDsRxJ9kVU3+iuGIdDsiALN80aoUO0BhDUPJEQ+MmVjgtzwKHHpDoTBnBFahTOMwXYs9w
sFHMi3FSSHnxByhDhuQU9g7HDg15Rv/FZXQEtvmhq1YYZl4nj8sECZ6hnqHbTTb4sHIHMwpkuVX6
WLWhPqwhqKN0YYb6OQASi+4fIE4iKyOZaWRWia01/iHkhBvPhbTr8c2QXMST+cR1veQ0hJwRAJUj
sSh4UeeLJOEIhQP+4Oc1sShBXJ1a74f7asIzRItQGNppzTom2pmA8EEcY7AGYv6UiDUruHpmI4c7
JvNi323na6zermC1ZOsX0FDrOjsvqUbfDkzGguWzebX4ln5iu3/sTYAGX3IneFU9riFfHTsiN90V
gIr+SHuEaC0VLCBX7VvscqQltgLWaD5QD3AeJ2WdCDJ/ckModcAn5jzZ7Ilad7H6WkLJlKpxWxfm
kpybpW5pj7NDGU6oApXSv84sENF6TWhyT3BkLwU/792jDtirIMFcP8MIIwEacYWeDam08rqOKi+i
beS6Wo3tY/BZ03behO7Nq8jNmR5FslFCi8VFW3/MCTx1bNJoieqmNvgVrNy7PpmLAebmjZsnIZ6V
t2lWcY4DT93eyVo4aFuExgNdKCqipxZzsqCQib0dhgHzFplnDdBNB44/i5mfItfjWw+rWFFoYR5A
chOWNwEHkKzB3ivCbiPN9ISic9LhB2aofeOMQ/6+oeeB3SSZXpHxpRkK0Vhib5E6p+IUg+Oq52z+
qhBy0ftKLxE7rV/UT2lDfYzgyh7dd/cRck/jHcwZnKBnd/2xXKCcFjbF0veP6HqDh8i5mwbctXWl
2Z+nIjAFtuwCTSymfSI/wq3L89kZwsCor3NLF1oZXd900nZZeKfaF7l4cJ05FEEI4BkQLAFfu4o6
7kfL70g0pdaMFlW/57RbZ+Zi76HBtRH0t5WTU2RN5QyYSfit621S02ze44SMlSF5OehJMYGXYq24
1L6NbNUNxXAb6F8SQPiCoaETjnV5BrwJILSTdyaacftQkWMf9UfjKLerlJYMelrSaCLVgmeaHWCn
r/09uJwObmYTInV1zBDgCVScLE2jsAgReVPHZv5s14D+eS+CUS4cDnVJn+tBMkENK++NDwf0steb
t7NthqJThrCva89m9ysHDzd0nuIntWAU1WJ04sG38FKcSv97xN+NpV3GbvNckUehZu9FnLDiAGDH
Oj8QqOI3k6vRb4e7UMQdOyNrBMd8WHcfbsqYdfu5Im14MjaanhUH6SVZ9Yh2qEf8HmF6Ru27LB1E
ccUyFsk5LZKe84EWytn3bQdCqaJJU92fNV8p1hAse+hvkDq6fd6tlnFWyS4m8Quv3ttAOL1R9Zvf
f1gkkpW3WaNg1114zsOgA/pGSRHOfgTNKheIJuPpH6mTx3tOS6c1LPjaTwGZBbLSB8msRqyFZmqY
IGeTibqzI2it5Jnej8nB3Nuf6XHb/2EiPRXUOZLYX0XIt7ikDHjEXbmhO0j3KfKvxbloZn6i5Xiv
Ew4oP84toHnAAXwQ1hTgtT3rJUKjJfS/T84erdj+tlFmd808rKopGNlOhkCtfOE/ipxpTlA8eoeC
pnDFLfUpfjDw12QyyNmhqzdE4ieIUb8ZJCLTEu+3N0KupcHmO1pijb5yeI7+rqdZgyV+NHrfCApi
RoVe32RJiezv2TsAnJBVtyi/VUmVJr0OLF7c9MvD/Crqw7UDSsT7j7r5hEjna+0/AMfsBfdn90mr
6ziFm/70poVgbsYSZ6he4mwnfxlw6Fz6/owEtlEXALIs1XIWkkTg6uf6UmIsJA9MtFRAsIq0c/a5
oh5xchPRG19SHJhiYx9cexEo4vRsg1cZm5I6zmTHAI3JByi+7kePOkEgtLEEpoxAn/rPmp3Qt793
4c/KTKi7oZRwpGXruqnA0yELVkTsV+92WLRqrHHn4G/HEqFr/PBmeOcg44p/7ko2is7fAYDFp/o2
gnQqj9+HpNq+cxbHdEXrRi8UgPzyDeJvnPSZx+UK+nlOtiBbSb+tfPZTKvFRbkmqF5hgedkAkJwL
5M4vsFqewYDu/p3Pbu+Tw5NDNNj1XS7Mz4ppmkfoSGB7AMtW47tnDWashYDXvgfbVjYIEXsqrj32
VleyXXMEqJmFZD7TqrMtbSPyHthqgSyb6OyQqXlwHChqvdG6kCzB4s3hXVFKZHsQAMVM3NrAd4io
Ny+GUTI5cR2xPcKR1IDgjZ5Uri6RTtJNl0oVI3HppWgQVcZjuJb+8fJ5OxXfG9eKEzRKsQUqL04C
Jm4Ylxb614DDTRqt8TC9IbRM7VoyBVUtzva/z3RSFq2iRVGFpiU4mkrtgsMdbNYW9lcvP//yPXl3
6lqAtbzDzkAeFW0QKpjC4NZffRloyrvfwNjxdhL8YJSmfSIN8yPJsAt9DI6D5INWMa8W3sEs3PjR
UOJWfnVbfXvSflaIs5bLFS3K3D4CeE64nUaKbt85++ulCiaheyXoQOzsnUIXsIcUqKW4K4Rpnbht
4PpMJPUxJ+ze1VLhCmSBLUAC4Ubf7RBnzctqKpMX0NT81QPMN6RTUct9MXq/PP6vyuUXi26g244H
AcTHWhzvr1r+RxXUjqPOgekuAMS9uGRW9tJ3MQirdLG65gHwfEJSDVuoT+jrwgVK8lPivhobR3qr
3GgKmDy61v+QW0igh+pPfLVtfrgE019aKEoFcz5zFSMoCTPR1YlTPRzaKJUCsjHa0Q9H8wPeV42D
D1d8Zpz2Xu/eDjB5JJir4Q2Hom0ztX2v9gpPvN3XUJFmRgyv3V4Lcgy31hDwJ56gvp9zATMqZ2nl
eATRHq3IYss1DT7xepvGUQFFpxGDEnqG8UVu8M8r2WZkTcHAMDzpg4RCGqI+N7f3cpxMKIrt2RuW
9pfhB+rtcgvH6heT8gs3C0GwB6+NewCF0ecyU3N2ldiS6EYZnAynNcYbcs3wnvgBm0vgNpbC3eIe
0r0mhRagaogpG/F4Sycj2GtCf6+dYwjRkVVs6agssrVYAyGUnX33nBSi94uabMDBTe1qqEvtXsPW
g+ydT49UM4JTe3v6OGo+nl8CqZGZ1SgNlp3nkgAzvtIiB3AMM+BgWBox6bcwj7jCLYUOzhpb5Lsr
LOZKsevCJITUeK2kmtPw8ZdOIsSt14vC1lDCQNFdk57thINOWYggOqgZ75qIqBwG+b4nvVYejPqz
5nYuMnz3C5UuoMidIyfdVhUozU4MXVaZHTjH8H+tvuqUyhGgJ/Law5eXVFOYYOKVHSVIvaQCnOq6
A9sj+ObBZpy3T987OrpG1j/Ga9P6cd6IlfWyCI2dkTvRM6k21d4QGJPod52RGVl2t4XIauz+EM0L
SzT3Xdz5xplN0+d4LsXjb1nRI6XmvDBLrL5ktwMqH5/DKoVXPMNju4UkfBmsNzf1NQpbPecxMtXk
NPz1MVR3LZ7plHzCxqKAYpYbZgnweULB/bUkF/iDTohwQt+xSVlbEaE3WnriUIOeY1nXlmqRRlmD
fEOsJPQdFvIYjKGChT51BuzgTBXPuY3B27k4rv2z/n/FItypWgvDwzYlQzV4Jpuos3RI6hgMSSPc
RNCpNzpnpGbqoxiikpOCLrXcP5O9GKFR8JwQpbi5QOePXJ7jinONibvPH2byhMe3M71Wsr/Hr5yp
ME/fniPvdLsQl25MZhbY6kTup/4Sc24ENKJFzhIaukduLn/OEs8gc3ArCjESVDMLS832jYuZcCdc
6JyQEfT3rSov154Ias+y1a5rlaYkNpfGYXqvyokKItgR84z1L/xWyQP/9xb+U1OLJec/G9tfB4uf
ZtSTOsUyHUdgH9ifEVRiTv4p1ZiqDih/9/e30zUGJNZWCi7DJdlo/sq5xQ51HMb7LByHwFxtdwu5
Ui27gSbrg7lHscw4x0wedCA06F7bYfROqCJizIGJJd9BIorZzrfgEE4Rdc33cyvQmLagAsKo8NeS
afIv1yckgd0UExzKYwzYi8kr9iF1d4shjKWcSDj51HtiXxtvSy+0jDm3F6pUbE2KCkWBvtrGqKiG
06YYd/lv77DBEsM3IPnCdUT3NJKXNa/qT6sJmGB8MA6hJCYW+75DplpnY8N7ikhzrwTLJWUywUun
QiUNHnB+itr6FXyNroU7wxxCQx4dkHCAsCzezfrzk+e0sHd8QhHRdw6JFIObZywILaYDMXq9edK1
duvU1oDOUHI44Xrc/hoFMkIqUjYlkjRj4so44InLVTeeK0NmyvH2KNaZovIppIOX9C164EF3Z6nT
VvXRXxh6hOzYDtjMwmLUNzh+eGPSEnIULfNjs/VjooKOgszaW4bH+F1Dh1GdEx95rAz8+4XyN01e
Swk+i72Oz9AWgcMs/2Ito7/0Pz3HNUuNlKrX2r+hsHoeEjhgx1L6RCU7HTFE8kr7Td7tbfiS/Mer
sjJrr+IpKWzG3rSmKUNSwDFKNA3eqOC8WhiJiXC4amOc8WqUB7g2bnt7WJsEWiZGAu/D+AUuzPcu
Iw4LerFTjd6r1++DO7iwMkVoieoaPjR4DK1Ti1ncz+M3OKBftZUilYMLNRVZ5n6W2FpbrsHaQsSD
vi7UBN2DIBAPF9wft8/K0wERXrEvrl6CdrYxRbOxGdMZyS+2F3X+YRyVulY+KIf1LpB5HBjzRaIm
12/cTtrCykqFmDhzu5M771BfKatQ2u8caWRnK4d2zCCpCnhH/jjR7AI+5GsTP26mzyA/KfQ23tYD
inDC12W4N+3sXQ+zFZdnSmmes1jZuiV+EZvC9qne1cgvBWmZqLYyhZ28TTCrvvihSqG5IwEK7Jvo
uQrXW1tw8Depr3nWpiNGslvyRbCxi9uSh9w57DjZ0cGuBpNRKxvlswsYNyksor5/cs7GI/Er33TJ
Lq1qS86rPBpVG6l5Tv2alyZRTKS9Szl/PQ/EM3loZMB2ZLKG1IpKJv/K3nOdc4o5GQT5VYmJgv+c
f6X5/0VH7MIR26gO+gBYs5kof/ucbzbhYo81b150xgO520ZIqmqbKlZVILgYJ7A2uIFxYCOydL4p
h19FTdHBDKJaQF/3rMxqAWbWjdLRt8FEvrMi/DVl4EDoMLVEHO94rs6uQMWfBuQFN+ECyWyoHPPG
kzcNFAhM+gQ57MBfrEcmNkbQ3xWiyYIOos7sC22IJNcR38+8FbjoKxtAQGKYhDrBDTAdrEOaNZ9J
3kQ0WangQlH7whfN1I5UTrMmfk63HK0ackkc04h8QQIpoz6g+Sf/7TvJI+WbLCVvJ2bFADHFQ9Z7
mN2FFtfYRyVIoDEMnl8hAIk5ylsnOFLuvMxJT3IiO1ee2UyCPlun+zIfDBHEBbIxentGCg9Uv7/s
cnyIvnaJCQJetzuHi2CcER4tl3LJTiuAN+Ml412z2Kt9Ur1/SY3RZL57pXbmEje4TOZ5m/+uuwht
i+ON0sC4UzaL3hH0mwhWiN4Rbt9ZXGS2xQZ04BoM5z9YIi4Ej2sAeOpcxqq3TF3CHupF+Ystph8H
9Jq3h67Ca8lsi/X5kfjXjdTBgHt5rwJowLyDI2l7tulWd0JR8XChRwVJoR4n9zd/yqVl5R54n9rk
e08Rscpjupb1jeU6yPY4mM35plutrSpndX2hrxsgWc757IMLLZ+unL9qYSZXb6B0hwSK5N9ODLi7
vTozW//4uhqFj0ddSept/PPE1jMDnNwTHEjidNl743v6KC6hRh2cMUgF45AJK25U8Pew/IijnHtG
G7NPQ1F/LB6W0Gk+r4dYNIqK1U0u5/seyqtYnH+E3+kmkNcb4U0goazFcxR3ZxhMCQRIeQu18WKE
wVUgj0P/Ozyq8u29wYZKKDSw9e4NjfuonFfACpVOCxPAhkmsKTVe1+aoaKwuQl8YHluQk83zYQo9
7vf1DtSDiHZFTG+q9Rofk8w1lLbHw8n7FcBOOi0OOYW3UcCpNqHk0yhXaaZJgYgVXgsnueArlQsn
eMa2EbRzrCZrRGqdyiqYj9CSfTB9wu3n1HHMGfIG4HwOBAOoG4UfHYIhshO1iKdjZXhRi2+KIGQQ
oRiiQy28stgG3b7R4Eowm46mpR7JO2Y0tDfR8WIY0iQnMaMVdiTqVJTfqSHgPKm21viTqLh/WC56
+KgYiGQlS45UmGuOYVvQ1OYrn89M8ME8VZcfJ52xeZgI1Tpphe62+8J/1D1JRaQ/dUcO9ybTarNj
ZVWO65jmuHoXf9JMPbD+arwb5wxAxcpawVMEiY78R4/8bO+rWZwzCXwF84LRNemJY5VQL/huKFpV
omTcbai+6fuKrkX7DLsrNmw0nu9b1me2m2Pcs8aDCN4Ajrg+K58HMIU4bNO/GJltWA2mljuIKl0m
BzvyK1snOVDqnIxs+gTGaybdcz6YNKq5J3G1MBh6Sw4CrrhKhO4gf/MDxMW+9DoHSiSJNGw2gFby
ilNgtf7AxOQ8mDKYjOBt3//VU9Z7s05TSad6iyx+xumVsrP80Q691L6ZQ5/X0BvES+7YtituyFAE
W0+YQdN1sLmq6gh0sYZP7rBVLuc6/GVgSJhD69EKXpch/WoxeZ2FNMe43yl3j6mq2mRuw7QGK0WZ
q6iUN1wK8uwkARW4XUSeG76YsXLfiOap1DvXz9AbMozC0oIi2ex7KY/bDuT3Yxr6y8G70BXbpxJC
tlnvjEd7nyqPdgTcG61/CG2zXvgHMLmnuqdoMLmveSrxwFjjbNFfDrD/UjT5n6Jpgs/e+wi1Uvyw
Wu4+pdmMB07BIxdiBfpgZ0Rz2q/NvqogvVoPuK7GfLy1dyAr1fF0QKhBLKpsb0eRb4wytaC/nMSV
ZZjYcIGLFHtls3W4hKze+aPZr0Io9mnPBJa1tuSEB+S/c5fhzH8odzuQMps4gNq6PCcvd7wAHTmS
qQgEjokcXJU7uMA0tARLDOqD8ECiOEN6U0iDD+cCnK+J036SQWPdlW+s+hDUlJ0Zd7/qU1FjZpWQ
GKtBuqq97/Ar3rRn2fGIqv7QIR106Tles3nIxgDRQxufJ7oTwKPYQa596JauvLVNSw6GPCLh3A9C
eaT/PF5mi0oybgnpB1cJ0sgk5qSEMe3gElAJpkSsUZfdHubQfukD909Wo64cuJTKQdYFZ4BXsxGf
rZbsmAJAk8gYMKvXpiOgZHjnphSL4BdPii5bVa59y4rjWn1pees3ZX6JnyYcNZxTff3XMh3vSK8h
XiDMyrYaLwuChasA89qoRjo2gDpZyLW3mQQhhKLnujsLaaaczjWmfvb14sE/tFg12Z0yP9uofcsb
g+725JlPyv5YaHP+k34GTIi5BHKji7ATzrchILxP+nx7zKkCZq4bq1w30KneXNIxK2LfhHtScgFB
8Z++vXs+ai1/S3OHu2ETtw6rkGYy00LhNCMPPY5ipB7WIotDqVpORtM29kK8wOBA/ja77fgjsNcn
DC58wSRnBoiqtVwXXTsY6IVfdFm0FHIYJIv6+WkcEkt7SSj4qR/Cms5KnkEaqkKpa3w8FbcJVGPy
6nJBPuI82wVnc/nMHzkDSq5S36HTcTlE1yW00BBsxgJzs5kfMjkl+2MWZqRpfxyugVMNbLgBnsZ0
Dkei/v3qi7XxFeV4mHft6huhRvyUhTFnYg4GHS5mCpn5mSIGqcFJ6VfAhyPdcJ2qr/nll+L+NfKX
zxos6tYtUQO5+DuqQvQ+FQUySy2UbQ+NaY+Mz3tVCuPOsmVgcHd7GOPy48jEn3XwG4SCJt3nrxJO
jxT74CFK2uAxb+kcv7M0HZ0twp4hlmgqkuTe3mAtgOkm+QXluYvTHFhOE4JMleIU7PIfwBWBk1/6
eBDapPuTDtxfedlm8gtjHhe3kt7Y6HmgLyoU1t5KQoeFbwZ25+IDMV7u7vb6+0bMejF3tRdyrxNb
a9s6hvUQaUQOQreXN1rg2H9/p1HlwA60CHvO18qbnZJn7Tt47mqUkLdoEPVxepcSmeDyBxFiHAM4
DpmQ1+ymz/Z0SBTFbq5GPVrE3YYJt/2WFWOwz0rZM1UAhWfk05kU/m+9/4b/hxw68rMrT5X67Trg
cpPcLRSH0SH7dpni2uKalvEMNmPFKAJqH2zH9mOLFpRG881PZRcPltinhr6Vb2Ct+6YYb+FdfFqf
Z41/x99UI/4OnoB+ODIJ0J5YDQDJqnhvBUj4iwJAxUnmZVrH92NVa3JVlr4ZMWc56VO+OFipjCXH
JiI5Eyb+PW5Q0ciQv3lpl9fjwjlZ6xbQN0CT0WsIACbgU7WlcQckG6aFK6CefNgLcZOup5egHd/K
RQI5wiMaUNOh7DN2YSRUCHdR/74YUpgNWKtauMolZ7XRPFIZkzRHIkU26Iu2D+/Ri2qFXNAXmlsh
EkpUyl+nhlWmuTOfi+r2VJ0ZFeH8QKbAuNKDzYzYVXyt7vjFgFJ0v5hDzTOgu5Q0me5lUH/Vadua
j831pNGOPB/MtXE5P457FWgWyjUAlI/RyGx6dvuxrzZZvf1n/gHfcAb0/leqjb3O6hrAkpeklxm1
GFOtr29Lf2HkY4983MpG13A6tvjeu4LgJQAahCVfq/cLUG4NoPirkDRil0YDKKbOx+BhFYTi8d25
4b7tKHZPZjcFaacTjx7Nrf9Daz/CUKXBqj7kfSv2eOtWQD7Oexv+wQ5T/8AxDUF0hxNTzdbeZp8K
QUn9Kh9IzW1WdvQcpnqfdU9FFhYIjfTLdxKGqckUW5NvKHBXoOjikbyfEoljW8S5p2y3z705UyxV
pYtuj/jCgWeI2oH7JzY7anj8zoMaPMiGAaVcDS2wbV8n1V6qFb7Utjk9h3azS94OWuvnSVoiDexZ
gxWAc2evgnypwduJ7JqHU8KYn9J7DhvzSDHqVvypLJoZ310tGSSl7WXMdpskG3Su6gcgPLuhZzUK
QfB6OYIOweCWM8+FRoPvBQWSHd2xzxaA+u2ba9bkYGjQJa7l2jKDfQgFnL167lBJmBKiLlNDnsMv
OqdQWNsNVOxxCGqht1IKRy2nEtbQhys+TA4kUjPUlY6Cg1XpAEXR/FqIXFOudqysfzmsiMQuZFGZ
Ejn5gUMkktwnTJCUbutLy78PDH2XaaUxeZw/gF17+wjkLRLzlcpr9YGHEgiksdiqOPwpdZXjisV1
xoc7UZZNi85uDxDoJL2TP3tfdlOe6lsUqWC7ZP9YM21DD3ddZayDpUbMjaDSqM/zMlYP7Dk8WmXk
PtWGQTU7uA5N3y2bRCU1S6pslAyx1jtKtC9PHYI7ujv1fEu4oQiL1cWEPfcbDu3foFjdFT5ABybx
Ouw2XLjPEHKjAZxtk4ge3u48zy0rOG5R1bz07gVYMTGS9YAtLaz/iAclCx9woJ3EWKex8SIalL6M
McDq+AIntLwB9PyxhS0XzHv0t1mznVxTVwIJ4SHG1BdETbA2P9l1ECi/s/ktjDh6q33R6DmcZmtc
oBeaGw40SkuccdIKMwgB1y6uUCIPxn4fSedPHor7PIDHPnAsk71kh2mwHR98/JkrD5y2d0HXkh9q
rWwutHYlAgn1kA18SXns+cmWu0TRsrwhfcBmqrfhQAQai86gJe8aqistqTMZFHFjxNo7u0aZv+FN
zdo0WvPlWKE0rwzEvQ5g+3wJlJvfXCEW9omabEXi2rWWArXfHz1syBHmdQM5LrU6pVdaL7+hvH0e
/Au5D3Lkxxjuir7r/eXSWzQHySJgaV3IgW+oMoB3wFuD/NeKe8ssCLEUq/0NiNC6/s2fE2r+fuse
H2FpyRzpcoSfr6BETQh3XYRiNWpxWqqhECZBEeBxiyLEzKIo5tFJ0gDR73N7fYJ+T+swSpuYZeVK
pIbm7WnhF0zxoLAPwnW79LPqJBw+MOEwVS0rMUsLCZtS+wyBxe+u13F7AvH9MNVHu9+WU061Fyqb
49vgsXmJwfG0/zSeuRWe3PruhqmsuATDXCxfWjVoj2/Gi/+vqKFJeFnTHmgz/zIAH5TBJOc+9PUz
kUBD7ib1dYI0cIfnWXbqfVBvIy/knq0EEeHqi0a7z5UQnEfYabmIFhoGDTfxrf/3A4CGA50Mas7Z
yFbCcKudoixbAO4GBXyiQx9wmRr5P5Jn8vvJP41K0SckuCWkX5FFZGFe7Hf9xkbR1NIblsgMIUAx
dVdUArGT5WctpdocWgcOIFe28AwV7WyLgeL7JzOcLKliIIfm+xlSj04xRrffgrKlXfjQIEtthtHR
Ee7Dt8HAkCvW++PER/Fxx8HyuZ11c2Jv3m0ke7ThKahwSGWkoOzXax07aQWfXr3swkoZWqhzL0v3
btC91buck+4qmnqRIJyNExkdHfn5EbQq3DhZltU2vMA1HuGhiYSi/nCVZjSUZ1zE5mENClaKHZvA
hlHwNMb+KtHgDLGcRjesd2Yl+NDMResyTlgbPIk1p0lWKDWFlm+RP6ao6kJO2dRDKp/d3AoC7V0R
V+TIcLwDBgqCs89LmfSA7x44cjf4a+d2J5FTMCEbAZlcQJMLwn5xQ4IBkyQxlf4hHqv5qPCmac4k
5R6a89jbjXNC1Vrh43S3jP8wjxBhjSVQGLPuG2haq/bN7WLx6iaMpkojVFaKhAXewXUqX2A+2UXM
6ORVGohMDFrQH579cOvtlWlDEiyAAU3e6F28QwSinArRQ3zpe0Arv1Xbv+1QPgstWtp794IIGDIR
zuJNmJzs5S034N18nX4sr795nr9aYrJDICsnmOSffV2XUV6ZtdgtUWLRFqZFBmnt+/aJ7q9AutU4
JtzKtq2miMDMfyK1suLKkB4jRK8lkjR2ACX0+cDMngG4dZO6MLiQxgbyk5MMfSsg4gqO+bs415dz
z4O6ONBR/izmK4ZRjZIP1a7KmaD0vMS4OgwImqZux9FrWK/QrDTq1cfybZNKb4tx4rWzj9kCeug0
dOYKHpUNAGLTx6MFvfEh3udq38RYtiZ+AeuE4NPVZjtkXpFr0o1lpMaf/ukXFr6hthVASmKJ48Po
SwMnxLO3ndu4WWwhYm2iJh/ImzE+0mrETN/hZi2siPLB2stgs8f0Tti3BIs+7WykcFcgdf9gK0Lh
uDE3jgRv5JQmK+eDlMTMZ+d837+lZxEa8mRZf6rpJEq0LIP9u4UOSixWQeGP3dsZeenL3IclW1cN
4KzWGZ2ZThY2z5KHdAhvYuOhJSZnZs3q5vDkTwxLjgpMEHUpVhvpPGHl2dyXZ30zMUQfWtFcoISP
dEifjX9nJCRDbmyjqx9qPLAA1S4L45Lubfi9NLFMQXryrQLMQJqu+7GcHgdQk7M34j0tJ15KLgvC
819e9ZJ1uR0C4p5a2gCOQNEy0gYINeMjINOrth/Qe9+uriCOc3layLuY8zgablHav8cg6j14v9Mi
aNrLmtO5jrWZdtRV1xQbgabh/u70hAAwpLOPCwHz/M3ITKw6nC4mLTEsQySZzkHk9mIpC2IJY32h
mtS0uUx4MbMHG3hhU1OKey+aQ42jhqEuz/5GawNZb8b5WSSxgl6q0Mt+qCZLIpGvvpgCyp3S8lEJ
UDL3LmNHpWEKOJCuNsVZFZ1OpWjEaTYVGQOHidmGmHxG5ZzMkP6w5o/7LDf5cQ/CA7TVdzVzTzN0
LD9NB9IIY7nhgiQcOHF+Z4SHQwSO135aInwyvQZCDyMh+rEjKgbHpLR6AXC7SbWc0Tl1KnB+5xnJ
DbeJdt9nr3ebtHlR8Va02SXuuDCKsWcFTSMppk0RGqieFZTCWd51ot2iEvLlv8FAt6kd8RfOyrIA
7mTPQwTlNVANcfpfPlbBc3WHh6aEnHeVuynP460gRxGGlp2yEISGjp5OsTloVuf467u67k2hd9sO
6/eZSA+OnYZVyMpMYrpblBpxl+ZzfG/sDHtlO1Choyr/hO/x16hN3xDYEtkbZVKGS/4z9DzXzJrL
TRh6eZ4o2kAY0KEC23DWa1cAJNyApQoNOI20eFTkIHdrAl7sicN/7XO6Q/TgT3yCY4gXNlLyGM/L
WTVGxhzHM5vB1kCwexvbxZdFu9xC7q+JdEOrswgyRWZCBZ38WwBs6bCFTtVyiy+La+J05wkTfa6m
7mZqporKhITvBmGZ+UIRfV8BgsvMq4eIdSCwUruE3hYG1byEZenK1epk1y8vtGQUYYUJeH2OxDyH
OqwVZt4HBoSrBlBHqenXQZf5aQ6wz0OoC1SkVR3VwUYeGKw/znw5JGuDz0+qhUYURnmFCRzKdZSK
6qFVy9LhfhSQagzkaTAtugsr7fG30nTpDLA5nsFV8B2CT3U4fQNnDXAG737METvwL5YyHZGfpKHe
iI6ktpGuQO6xVCt4xfF01pkjrJFaDdQlwmRs+K9W0CKKZKhH8SY/U7RqlpKBeRTzi+rFzSJWwLQu
yC6Wkr7ZOxvnpBhX2LAjW6lB2MQx1qFk44noTmAWeb0M++yW004oRJkpqIFTuZCAONKls88Pge8x
prHVTxVPQXuU9UMOPDcYyAfWRv/xqraHLIsp50FnzNbOyb4jKy6MrQKyt8z9TiBiVHCboTXOtvlc
YZht8R97v6KYkgQ49RmwmRq6urHLAVOpWG46u0a3b4AP4Y8VYbXN1Snfp/xVYCxIUvBsVjyRDvqO
OvRlLmCglSE6HpNP1iEi4yayp6CuCSjweIYA+T7swyHKfGEPSnDvUucIU1qFl9NxNQ611er+ANJ2
lCmu6zKrMd8598KNDCto7YH3hOf1r8RjoYQX+L8YrLY29c06rbt8S7J6UaT1oRdWheFOhDZvDqGc
btRsDGr5BAh5zXjsXfEZ+T/u8iK/X5VqTz+6vcJnA765dYPacsgWF3QpTTMDy/r+JMpx0yUzWrR4
3+F///Y2pz3+4knPXHCHPiaR6b+bCaZLkBv/48fWimMvQ9zQAbQZH7cvqLgrKJzm2Gi8gLRTG++G
R74x1v3V9eUIPteGxpnZ/idPfrfk3rpDjd0sn8nQcq3/K22NWEREw1+eL/LpX410R3eMjCPm5Qe1
MX86MMVFRhrScEmreZ2HYLzH4Zs9i78Bm83gHD3xyvMOHg9NSyroIW/Pspmn4cUfHrwvBhMNiz1s
3+eFCwXiJMbta31p8o026AlWNPlPPQzWUGw9Mk1GhZJdpmgUh829c5+LY9uFcenD02h2qBCkxrxL
TI7uL1xegj9e/pjdSnoxQNXDXlcIPH9ZQZbAEo60RGIqj5/B11lXVfT1r0ztDvj9yeN5npjGpSZo
pfhcDSpAH96DZzfQ7Bgs4WM2rzHTK0KweENBb8B19zsSQUKUyO1msCes0WIkaVFMbj4N/Tb0XigB
yubx1nhwO37qFXRDbSTkdevHbuuXIc0l3LqQnwN97SoVSJfqlF3n2BJlKCaLEDsJNczmMKSLABWv
X2A0E+ryIsxKq2pfzn0svP1JcMqrNwr/W1xe3EiZlsyIkwPCnPnoC0sJNCBZ+OeD0GR0ywYUjxDO
RNr1aJ85vzh+JKWYpfyXDESJLgKYShHMet3vfE/pUhg3XKyzry2FH3nRa86+oRGZvcvLrlEjoM0d
htteZUyLZMIN5w7WTYxhyYj1EEwhwPSbltPSmrIjSk/nYPFLSPUDBpThfIjKRnRzEmXfAdbiWtf+
cEzlTO5mBkbZ1J++O3rrhXgzYJ/e9Y1PeW2JWf8BWa2gVuPQfaNRb3m4iXd0/nwpwFQ5LTV0JqaL
JM5RJnOKQyLwg7YdurUh3J3UXYmJIsJmDa/H8Kohiqq5QbL/h003fdVBRlDLUvnTpNPN5CCfH0z8
7pV59OptSG5Ox+2f4BBgmiGN0mW0jGyBvNPf8e11n+HAPM+fo9JEubsocKauA8qaPwixkA3CTi3j
MoebHksnVjXTsWYqVPkBACRy6gbZvOztAbzpiiQ2Ctbeiz0MNfnvGxPWxkyCl16IiNv4vSrhW/At
2PX2rwtj5GXmoVAli+oyS0vAKwHSp0eqq5vR5WYLqhM9bXdnE6n+RcQCXuYlr7R1H/myvSpSz5IX
kzMnzUlWS98UZZKrxGAXpQH+5ddrA5mg5yicE5CPYVy+7i+7sq0ZQJlGnDtHr8a6yTAf5RkcRZON
sXSt26SsAD5TutoCki2uIcEuXMxgdWMkZqTgiKsb6dRlWflm2lj9q5aOnN/BxDYMgGE9Xgaw62My
kh2CP1IYa0L4JXeu8BkDlLDFVRI5XyObRLPvZPA5SH42Af/WGjoTbdwV79ezmd+IE9FMV4jsA5hZ
h7Kl3OwN1Agd01KFcVReBNUT9DquWSreEWnGpCDMyABi3PImRhITfNu+0nbwB8kBW0OQf2HTW64S
j9bIUB/6Mpy7ZRw4rkxXfzMpF/eW9gzWtD1P+Kz4c3Zv7WwT1RCprbqWYUgF5HOwFnjtjG9q03S0
Bpm+jLEyDdIK1Rppmu7vWQ4oJH1yhCSqN6bNm3HI6DPdjCkcfgQwxuSl7J1pnmjeaOC08oFUuBtW
NQLgsIOD121jTMQvJTafeZKhyM2CrowgTPo6U8j6JDOAWayjItBg1Y8jyBhysvRJDS6neziJ/7gu
ADo+V5JO0SdMvQ5NGyfxDJgWxGZJgZT+QjKJpukRqbIksc7KVcBXrDBkONMChWjtQIJkAknsBp6c
w6r23BScQdH1FAR4CPAreefLsixwRFQYXXwwD4gjlfk9v/VVGNaQ1vdGCnGg4PKMSYvKfPXuAqJ7
x2AF0AM4YvVxnFTx+E7hZlQAqWWBDL6fqMUDlG48GUp+pxY0N3l76NNTgldsSjQC2rV/fBSLNEpT
9CoZ9bprUQsHxklEB9Dp3NPfnVVJSdxJVl+xpCJhHhMjy25vuperhDE+xhdz+cZWgn5IyLv5I3L9
IUVGcS8JI9ZF+pHybRNq47sVnsHJHRRp7C1DWJFSHljX5x3vopjtKdwy2Ft8Wy0Kma9zOqZ29Jum
Rw6zyjiUSaXiidd2tDK7lCAK8imnfr10b3TJqHShBZKJBUx+I8hNVgK8M0tJm1jvWR0kxM/qmN08
pqT+vN+J5IwX4+h257MQSFMtzPM+N1RMqlS/NZs52z4dqvtG2uyUZIm2cx7emsPzIbeqrZIFs8PY
PW8X+mYV1V3eJoeADS8I+ls9ZcWVzq9BDBC3iztdTPruXbBAQYG9x19yYRDG7/WPZXBeWToA1mYs
c1LDfbaxu283lSiAWr3Nwm1+HXK6AsM4o1DryeAfwBt7zKldiopRsRVum+0DGMn5U1ou+KsBVumJ
r6Pe0DB8SyfL3hB8EaY4JJWDSoQaYSJY53nHaamuW/476QHDnl6ipfBi29dowpo6ww0Lr49o6n3q
4NDru0Atzfy8bwaYmMwgjhajq+tAZMy/r8oEI1supq8+HsTcHamjgtdr+o+wvFxi7aekEga7CAPy
M45D4rylkmahAfFNK05CzRS0wXHCyPIHYi04PF3H5edoK1uAHmG8iGjPVKjHh1vnvyCDdMpzFSoK
Z+frja/o0t0sbZ/Gg//HErxPrEDvoYQ8NaFXKCX5PuWeEps0JEpAbQYGFHuCkKsYKsNsZzMxR0qU
UVVPLh7fGUByyDnub/qtTH7q/oPVBpwNt0DK1gZKf0TzO1+PthGQrjTorZyyT+ihhUq4bA1MtX/X
0U4NRIT1wic7W/X/z9H31ptTW5q3ZuZ8jKR3OAKZwOy5rZeJ130A/WfgzrrlD74V0Q3dNg1ZKJiK
bNqCZwA3gef47ZvUSrI6szyC/giGL5sxhrRfBrihMhDzn4hgRQd2qHkpynAwYzkKOcLiB0C8Y0Hc
wseOrClOtZ377/+f3t28VMe9SIQ30bzWk5NKl9MI6uVTztu96NCgwpGM1CqplbVeUsc8LBuf/Xqf
J/UX8Y/qH2yZLF1/kGq5GsNtkiw5XDDBU+r1jOUio29FZvbGA5+H+7nxLtTUlsy7U7qkgAUp6eoD
kTKX+k4dcVnRdI440uFQl1A/YAOOLR9682s9uSuDsdsQTbm4XjVcil6AKTFlxhQRcuiFMrkY3SRL
Ll55FquwINhNkgqQJHWV1c1RAse5zeZpWeW+uABwNFlUZa8s9iaaVDmWY4ayQzNpBYilhoh/idYg
Jw2R5wGkkx0bq7s8XELjIdITaSE7HWmcRBio+Ku5JzkfFPxVMBvS1zdv2yyevVKhy0CmLHe3zjk0
4/fB54Iu7dIbf9jS0GX9EojaBA11bE4jmR2u4NupbdD9B+Jbm/mniIrTCscyDfNRZ2yQrhMi+A+p
hOY14DsekverHABCgWlqUS4jnfhwjsb+IwYYtrKf9PYC6umk/GhzvPcjiclne7K4Duz5uOmnbpVR
VkGsHjtaMWTppHpHrMrbgYK+6DnVLbpzl6Dg3tpbD2ntnFP9D67FvZpOnoxIiqg63+Ouy6SvY1cg
dvvbfilM+04goPo0T0Fmxk3oi2B9SfIsZ10IfEP4qSr+qc0YAi+NBQNSC3Dkak+7jOPthrSNK/Rh
dwLB2Y6+qt/+j3BCr48pJB7Txa/7JbO0TCVNQXql6k1aB+oYoqvclbHsc8ojyFCI+UvymL+iJ8d5
mFqLJVoz9VAq1jwJZo27lME5stnDoXOqIcEuJIP7BD7zlqvRZwrT1r+I+CS42WUomMQGNuEggSM5
pJUW7sbbP1rQDoN3VZC8CcTt5txrbSi/5T2piYcESL+wLBxEGn0vD2vazQIaCKo6+U6yiSnqrONJ
idGZGRXl0IfeZ3N9pJvdt1ZFdCYw+ICpb5Hw4kFvKI2ruf/i9nif3vOtL96+AeUxLpHvWVsY512J
0MlPh5WztXhJgDdoqsGXCrTXdvVydbXuwEeAAk1f6tZPUEkUOedQR6MSwBZPFTrxjDvJVAqCFRwG
XpukSqgFSh+kncg5Kznnl4hC9zK3AUDzVErv91ZmfLTmxCgWv/ixACP+AuMZVab3xXagd2DEi/1w
NtT0JkTZ/5ia7RlCuyQ+UtL4ZmqJu+xylYSX8Hha+p31zqLOvWxyRUkDSIalvGJyuJusjrhos42T
KDOXcapKK8KFTHi9PGoXVNAzSwWZcQPRqOEkevXVy7DHcQ/m5QIeCmEpTFY7JtIQ39N48+Tn+3O8
syMTun+rjP+Pxjv1OHxGU0gnzIIUYZ8lAPEmkKazXA+epxOeMicG0RLIisOiQ1QpAm5spcx5fxR/
ua4s6XfDBL/jyzF004ksHRX5YE5PMaJLjYU39XBdltNfBUu0Lbo/p8LmNYV4ywxnrTg4wesWLRzN
dP7LX2A6U2fdsorLLAOevEYoUSYFn43BUl+BTzzuji29+lCfHxvSy4seSuAX3kEDgPgzs/yUT7Rl
/ycyE0gHZdfVOkc3cFDK/4kxqlgR2nSOGFqI0w8aWkDTKsFOQANZOOWsdsH15Ek0Uk7mtjfAydYm
5qQOEHjKsZVCNLs70jatzEe2ngQym3Q/8x4eHHYQsYV20V0wqMS2wt5iSm5SOu3bTeLooPGLK7U4
FU2TcL5EWIcK6QcmVBx0ekNMGAVxO0d/cJHJ6ufMhxDTJ/WsZc3jJetiiW85ckjI6VE4/MuDIxbf
+Cx6F/A4o/6AL7z8Mxg/FN/5yAEsjq5YqMY+LWaaRnP4KMLM0QZGwjPkTD6FyqVLaAknF/gwK/3z
UNxlSzvjcZtXPY5FerD4AuoQ/h9Hs099G7Q8IpzWRcJ+HQW9ovdzXcwR9L6wMdLI+eqWREzRLIdm
jbFKdgrtwF425YjQB+LfrHg0jrTjnVmYZsBBi3OHdNcEqv0k+nhKLYQpWY9KLcSnZsAmVMptvugP
WG1abdRZ3UbuE+m/LD8KLD+b6C/Br+Zi+slmCw/3Jvest3wbusJlLyUoJpj3G8Q96q9j6WmJwvaT
A9vABqvxdy0XYhYPjJcmG/xvV66Y0yJnEMnDMo5dmcfOXq60nHV9tMPh3gHfZrYGBgSGknl/JBKV
kGkSh6k+Gehvy7zIrgGIpVht95vibpHWMgrbz8PLqTwxKAZmFNtLn3EGUNuyW2FISGv8/N1KY6XG
y26lpQ6wsRrg4uIPjmw8W/K8gTTs/cq7tQoeyr0STPEgsG/JSiGKsbSvympi6EJXfPcBLQtzxbGC
c0vOLPYxd9oZqMc48t/1CUOFOBHTcKxcXcyABHDf+28CIrv2w1C0wij1CsRi5v1dVGxWLh4FknuO
an/R/FwnyMyNnBQkW6sZIMEALr3LcfgKu6oGylb/d/zRkt4/J7bT/JUX6mfgGRYzk4CYZE5f72er
+0NBaaGJ6Q56wwVfOgvGL07PW9bNjeAuzAtmXY5Hxvo2F+W2baoduuqRpjjSZ9BkQwTO+Q6KR+FQ
lXOfqL7s4yLYJbmG0FvIMU6ndrIhZJyaCSL91yn3Tu9F4VZbSuXBfI71TI2Si2QzdL4FUYzIDVH/
SXFmEBwWSHFBF7wTef8B1Sm1Vn+8pJcK7CEkLLT5DM6kGrOwb6dgPbiR/+b6FMgpDhqYSVCmlI5w
Pa4lgj7rrVzQE0+UaeSUqIfFT2AG1FRJ3XkPWc1zj7C667xBVnnBHvcA/qwY0xxkzzwvu6uBJQnN
l0/DXZvPj4am1ySN0G0zkMJmgK4gQso1Yp7QkW3LAIb4qQQUnCGROA+1UOSsqAKTzIh6cOexNwN0
Ol/bj/VS0ntWgxZLfawMSi/e7j2wsHL1xLqzjdjmzq27Et85PwKscsRTSvMBQKTLn4GCzwKGiW8o
hFu/z06zQym0SI166+mGj4tTcfZ3sqYdIdwHO0HvbjGZEDolGupsEhI6cQOYm3L99tDJJ9PFgG7J
oUUTrWAeNnEO2q1JpPtzVYUYGMRQuIKOMyFK7XOy29RCwGEbLerUnWrxP7rCvmYBcoVokqkW5wEm
LMAp/p1+t+zeRnxIryTVIVou0lx8eapsdzi9vWfdIdRSJODnLyPLlKq+pyGFD528aI4ov+fT7WlU
Sej5DVdTcfmO5dnumVsZrvFXYML0SsH2hIlTivS3Zir1lS1HR5AReScJ1dCbHEwZOnJso43KVYYd
hNTkIgU+0tFAuTMWbXrc3WYVYW7+aEvdS1ZQcpyFWoWWYrIVfiToSEn6wD8lPsrig+OZ9WwkrEZc
PNnK+e5MDj4kRyM+bSWLSUOgr5pSBiYXSQ9nzOxEslkP2gM8A/fPOoKSWdvnUdTG1m7cf7sGHbSx
id8LsIF39a+eg2MIsnGHFccSpUC9oogEUAkG6ejXgkTbMYNAHbctMmvnrauB8YnJ6TJJ9hVn57UY
ttZuOhmmGxJBsXTb9v8J0MFBPNcjaT9vtDi3yRo8R2UEshtIm9qhjW8EcAo9Vt1tIObDa6gcauNs
PbvKx7GN9POP74PzBmOL6mEhm5sDmnfeZ5d9C1itZ4jSodN++eN16XxzOztQEUH0Z0CX+ORoHlOP
742t8YBXft7PYtNL252CDRfO+ICqcSJ6vVxobF9VhdEhGt2QcHqiYtGdDAoJnIX/tyi1u5geD1pR
wMsS82UxkFTxUZ9feFN2+A2CnDOMOOXon/O8gHdGkrxezl7tvFdMHTiK9v/jMysu7WNSRuXNbZCr
sd4tx+b5NiYwSTmCrhZvd72vwIZYUiSxZ0MmRJiCm0WaNrIhDIzEWke7nbxGs6sENFuvmbbeB128
atkoe4cNKqo1n40wNIwE+JmyUKU7/GUlxY38+bT89iMfb9m/+nLMSWYwHu5rCwGOrbU40UlSqMKt
qxvrzkf5zWSATYybsJTC3OSksWtN4IuA6Zu5+/2BRRraldJLu2hnc0F7AVkrDUVCHWKp+KvgLQNi
NpDZe70Ch+QqXcssHi1FoLVMSGQ+15nS2uwTx0D/B6yYlDeO4BLPm7XOL2OtsFrwX21JS133tmIs
ehciT7boNmWWcSu7kgR7MYX81UXlcF/5n4Bwaee2Gll0otlciffZTTUIda5ixkFI2tRBBR6Bp5RQ
KvKCvjQfQSOa4QQjU9tBVBdhnPOCzhQnD1Hb2mqUU+6gTCV27qW4duNeo5RlG9bpo4YDTvra5ZYR
H1+Z+r+l+f3nho1zhrxHoVNE68fluzn8eUrLTl21ifwO98XaeGNLAnfREwPx8mznnSH3ObWk2zM2
bh+F+nLLOhk0C47AOXnMw/La0xkRyZxWc7Py9RofSCb0pfTQeD9g045G4/MQKN2PHW34HcbrikKw
6TxImngR6vY5xNGDc9hKb2MtXO+/DEw7iJhRYE62dbJJVgfaNUy7wE74wAcT8zPNLh+II4KxC4I4
X9IIGWu0z0kUr3gvJUxZQVYBfXw5WzTvpEc0TmroTKv7mRcN37R3MReyCvWeEokWsk2qQU9Vd7s4
kLNmpKfgfRbeSZM0ElfNU6hOG5FaB+M9C44dOQFNja2v0oG3U4pJpPq4YGpULNfLYJdRMAIqSKv6
YrABs4Ua06gHrH83rVJ9lGwsCDEIuQHkIt71ACtf5CTI8f5iBgP/+GOi51Cd8C9hZLJQeLF29cej
KZBonDQkAP0tUDCruorx6xGi+OE2w8ojp6KUZh0lE8cOSzPJSsdp9cB49tqyK7P1WKGnum8p+UQ/
YsBqng0/B57hHb5h1MN5SRGNrTnt1BtQYfSKPW4C27IUVd6z4R87FkREkx+807Q7pZWVwoSBjMTi
27B6YVgx87YU0g1TOe84arbynvIze3E1jmaI8xvyGuYIa4j4XYnQk2pBUE0jCiF7Saf7hFjyR4Tp
HfvBuoqgPS8DgZ9M0Ckgeybe/bv0UsofT5FsnCOztr7D8vYLGbd1yLBNVgRUlt1M0Vz9ppFxHwzi
3ArCqzUaHYM+5j9zrSuchKuVbirpCNOVEzwa1qOPJApr5uP8+r7XQ9QsLjNGhDGWsHelW4W446xY
k4CdknMKmJVda4EkhFpDmyPkmpYZdGKu9x2bpUk8t2+XeqjwHL9LWW+n4JVdkdslqq3tKBlq1QHh
fzbnJO1TljYCZGeuNSD2kZHA50H+hxpFwHCoebZa3QQKVWKdvgbz5rVcP82uChcQrtN+zdGacHe2
1ep+18C+yW/orUjXN1ptsKyqBQT10bP1QV6raw/L+uRgHgaQXqyk8wrIztoyBwD2tapTkIbz+Lxy
mkZyOnqyGy6ZR8Ot95v5hmbeWRi1R/PWL5fr4raQSyoDb0kL9OqhhxgRr4Kh+tqP/2SXnWoXVkS1
61LahU/5H3AkGEfQVmyUqlogLTpHBv6oOVhSSDhk+25wsupYWtOE0IWV7R9iFY7Vrnf6gOhHlaGc
fbOm6Ls+dqtt7rJ7A3ESZUrNpnoHU0GG3XD31xpxtxNyf25wfUKhoq+IxfdI268Duei3KPf8nsVL
+Y/5DVtQyhhWqeLr/NkYSwThAj1P5i8L/KQYrh6Ce9mwerFf7CCY5lPATMc1ijF/ygZey8nFiw2G
ohvP5fnUIEzAaOCJ20lhgeb6q6rDTH19sC16jV5CIVV064O+wchD0tCFMeycIxpukHBKK67rC6kA
zL6TOCbS5T21a6xWajw1S2FQsy78w4jXzAZG09HQgRsA9T5fWHUU3wDHyCnGjlgIVzSUz8QdlI4L
LyZUho8ZWPAiEq//tjcdOrgNl1VCTywOMESdif+cgnAXeGqylyqPjOGHAMFqoaIEN9FjjMlkjUCC
8WR8hGgdZYO5gozRN87T0CT7r969kAkUAq0JyyaorxcriwtH+CXF6HP7XjkzO/jfWV6wi+cAZoKm
TSUntLK8+x4Q4HmS7F5c6XZROmLQjZ8Nyq003Q32CoHMWnzf5rLtGGabLTYhu27YC7tc1fmYtrtz
ujWgyCTMJZX04v/4XcuqS0zl5DcV3gjDRBfxnjJuBLeDewXlrSl3UpMXCE2AImfjYGmnAsxZUvmv
4RAACHhBPBYoixEZ5FzYEMUmByNoBI6awB6UeSjcNWGMDeF2mBSsqrMf4ebwJZwvwQ9gFjKvbHWS
VprVcyx33JnwwOhRXR6u37tt5IIuPpo99UaKwVgdQwVmS9RZy5PjdaaG3RIbznrvvrMC8DXohAVm
hHLMGte1z1qJD2YZUp0IRUxxVrdibvFdqyYWcW8u7b49AredSOTJQnrnzwf9mZZdoLh8hUi32jLi
P3SNqgQPc0rZXlHupkcXJ7VKZrkcVeM0eqE3aXRLniJJ0YAR2uNFwQvZ0qcmfBOoIjWTxFKtSVrL
mrkL5r4r2iCdOvNAEL8cEx3ONItx8ilsuqNd8NsQfSyxpZuVI2zVjQDaZAM+/p+9XSUBPeuTg+uL
UoD/n/5UzhrZ7jYBgPzc9bGsQ6Hx8fJQGeLYIoD9l3L9JO3L7kM/UsFfXX0psdx52oa2cwFuxL0F
EHVpyalRg1pKOyaKC7tmq0Sn6BPst2ityDEdUbt31WBsFar9MpEasWg7/4EtPoaznBVc3//FYeDH
UHgQFVC3RKyGEDS/OpeCH9fZgUGXit9LuNSjn4iaaKr8DlT7s/4iuzv86ZC3qUas0DZ3RZ/KYKEz
k+eyO4W89ro/pr6pG1ZU5QLx1TRDx6TredgvrltbunR6gV/R/wyJgzx1D0AVBdKwhG3TN3nKQTTN
6NpIuzmU1ad3oNXX5Sfk6dH0vtemWEyNaoQlbavxocSLuFQ8Js8xV4dbDzFB1JEmSRQ4GGS7U1Ie
KOyGOC7zd/u9rQey7fy8Ievtb4Evuan+FU1yc6sLzaUCJ3zsx/178WBC2ElQGTNXqJds1BopQCPh
e8kPPfOnPVHccraqSFV6Zfq/o6wRWPtzbYc+Z5w8j6y8c3Mf2wJd2Cuhi1ttouKN6WS9Iz6C7nMI
BIbJIy4zgqufmzbRTn33JguEYUCilw5X20TJY6TbtyuiEAId/OrTa6DyR+HROWH3fefW3R30cpD4
bJxOVuZTuPMdP8WQuttXznT6Qf+38/B/j3+db6GYOmqumLGurVD48x2EHtReQctdSEUp0gqtys97
TFuHCNOCHqfllwg/VWEb1HXTw2B72E1RM2PTWnQ5nKNmdiBd3BJDKrv0gX/fw7pm89dkBSiIjdOI
TcT1ARafCDlXV2oV/8guf34/SJLu1+loB9YqWatkxPcrzgNZ/PKsuQznbJ9kMhFzZM+mOM0u248n
LxmjRzw36Ok7NMhNOixcAEsl+rlUGJoi/tuen49gr5bkJTJA5ikpL60tvSNpvufWMrhToAH7m4cM
bJPARzrQzl9+BPo7sdmBzX6v6rSDvPPVKAvNiwRwl7EogYA74OAqpVojb9rZkkE7ikHPyBuggL65
Rg3PPR10yVD8DYUafccgZvrBMak/tzwDFBruh6S9/nLghlA4TMs7qTdujzwXKW6ky67hQ4ymwQ+Y
ilLI9GCnJcXtdFQtSFtvNAaUO4h2AO7WmmCPj3jn50GXq9hVch1/0ZK/+ncW/Oi4RJbBzBQ0fEDe
cAwV+O5GnZkk7aDt9qhJpqs+K61RVzf7cEj/KXp3FTtrgLC0M2Ss3DcfdUbr2LSAAeCMMOm1kF2Q
rEiY2bW+VqZF8SpeVmkyP+Y0yM0HowfTYMKzEvAXK8nz2vBfQztFGh9MEnxVv1vi4i3yX0aNoR76
zaVluvEfEG9XovwfjYFC2EAppDmGlpgRKV4itAH6yQh9TrsyjTwQDl0BRUxkFCwIv4c+eeAkRv+z
H4b7ct3EM6Jha/BwLKQ45VMIYtHEYSl6NrZmEnnfrb+bIBFigMJ0aLWdOKagiAh8SLY5keVTr2OJ
voCCx1VHViR4IXXP7WMSzYK87X3w/9qG1yFHwVzQWr7JMh8ijlT8g7UkTCA2WC8RsgA8hBHlWPIg
5T2NZpVKUHnJXZC5PTsgE5xj3tH5IIG1W/LESVhs98XUGTsT8B0dvpOfr2nvQg34Uzc2o73lj30i
7ceGdvnRXsysyk7QAP8L0O66wX2eTnXcTpy99ZTbgDdC3ED3GRovysMw4/YlIUNDijkCIPXrammn
7MPFqqR5UvFN1vT6ShZN0pQDLEMMopybvjheMaw+rjGFa3XZoINPtUmYydFOhSy3cGWP+U74iaEm
whc7B99Vr8HYkfK56w7woPlg9iJ/an80RoF/xqh+P1e3GR3X8UdaSOC8pbA+POwtYqukyookXfPq
gFeo02adambXit7XN9nmexj3T4ODtl8F5Vk2C59jCyQZYMczA9XYlQmc69c6VVBumdJ6q3PiBzMK
sXkyBUyIU/SA/FP0Es5gzA22NNFysFqMjsm2i5XKleMK1Bq2FMsVkGk9f7z5+NL6UPTKIrNp7OaA
AyNAJfSGiD3fhR9hYO+hX3tGARRxub49M4vaHy6q5t0RLc6/w6s8XzVsppxyT4PyqyJWQj90FikY
eo4rD2S477Bu3YL1R/kb/wGLtv2fFUX2gTnys75M1A8O2QgrAaEgaHLJmRUgVeb+o1S2RPnrnn+j
IgcQgbR6x2HCE7vLOe3D4J7NTITe5UgNDRN82Z7Fcz1Q7TjKHkSwbUnPYPOviufgxZVHPB2CMg7H
0Hi4m4AT0qzVckxGuyhLWGXYrYdAciO1a/YrTYaOP8jpl6OChFKcDeNHt/w0XF5Fme8HSjd44nnw
8tQesnfc3SKJKw7LeupjpfrNC2lmnM8WKL7fEXkkF/1czvNoMh7S/Gqy8eplY0QBTwE2FZl8E0hM
eiWA1OL+FoxFOFFAqSW3xpyIASKShZoGTAvEP8cLA+GxDDj4Jw5Yu2FfkOO2u3eNHM8iwmtISZqG
GXwE/7jmr8WPjthvcs7Yj7pY0KZOifOpirwAWwFWEit9Lknz99Y4zE9wrb26fmQq/coXvlov5DNm
jbDs4QHJXl/yrVuKSFYtQaLcXQ5Xmij7OMeFoBDxH22v022WV10KrFVHgWHtuOa4OdD4V8MXJXpn
LgojqeVNi1JrUJ/a133ySLeJEvjtSAKBpB/5MCI8vRyQEitwU+VP5MeXXz+PSWw2f81OOovROUG2
OmlOX47Q4cFZDoy2sTwWqaBWfvmudnekFCrzcVavg9nu/a6En86oOpSWUQA2Xi+0s+6D/yTa0qLh
MOR9yJB9Maf5XcQWDyBnaEGyl/B39PjsQM7ETbR+IGk4RCOhDkNMUcg77ymDM06+L5FYyfUFlOV4
XiLaKAtukVL1sFM8LleVdK+bnVQOkgb3jYwPy4FWQPdxPdO+y8i9YIDQ7nDUlv0CxrZiNta42zqU
p2q2YLF7ZZw+TUItL9oSfBWJQE8zT6f1PsSY/rLWuTF8GID26rI6EsXWxpFw1EHkbltzX+Ny5QAo
dXQYneqT8+HKuCV0FnJFoQES/14Vsqo4vQ6asRfrigQfK3X4qNLFONNiI4ntqgNpm7gvuZHSa19l
pCRM17++f1maAAVXTWI1TGjRgDUJrndK42XdCYawbwMDTxoJUZSo9hMqzPjwlMxSm1DG197omu/z
nkhQYFaov4vY5LwKv8RG1ejanakM7KWpXMcR/yu0harQFxHCRf9u/ii39kbbFxtvd6kWrwYjs1l5
Hn/AfxGtuGRZxdVAoeKJ9D/aVKV8UbCXa5PD6YW/KEWM5hx1mj39QTcciyHCpn68lvTLsGO1SN9/
zy7pdxgNJxlcGe0bzgKqsYrQIFwBIFeZUez//rbh6q+pXjvDqJCBfxDnyV2m+giw6DdfcAFj91Fs
BRa04TYcTfzG5n5bN9Uzl78lJCoGOgX3v9fiDH4wxQyKwdoWvtQRL3ruIDRl+mDLdW4qG9vFG8F7
b2GCyNh5rR/7mZj9c3EKtliW43bqNiCu7QY+7HGyEngHspPeld0R7fINxlasjleyf/UYKKmEmIEd
DQznE7Gfn3RO0Q77vnHuUSBAuo5c+aw0IG+a550/qLOQQ7JqDmBlpgzST9M3vipTB++HOqi5FXhL
q8MPAU8mllWnnZiVI4LuP3Wd81+OLuwOwNHblEi35oCpiirbrSKAGHcIOGDNcloL3/swGC/xIekX
6NfFIbRrbF/Q3JDw7feQDsHZXu11y13QZsoEPpqANBr8rOaltyYMq8tTqCMY1046U2mqdoL+0sr3
rmSNfVjkMsry5pEQUOS63zJzdF6cW7bNoYteGEfq1Fn+3qqfIpUp/nKyglzER/AYwrsGAx1ytqoX
Rm9tyoYJr20FkTpvVb9oy1G3jWKpS5Eu2PSG+v+ZciFJQy4meRpFNN1dNa+c+lwcLxz2ta7FpjdL
4Jg7JBa0ERO3AeVNXB5/V1JEtpZozs24F7OIGfOClFNoVq5YO6egHWbZhb7S3YLSOQ0JQHqcEHpq
p1YDDsYzm5Bfy5GatpaQgXsmewY3yRt0I+nNM6Vg9tVpMOrEX61OyY+aLGfHEZWBUgwwYcRMXW8d
G0Fyb58kdCnZk3Med+2BNfzJB7WXkqvVWRg7HipM7vg/3ZJ2PTrkzVb/p7mi0JmxFUIn+KeB3vkn
D02WeihCIQbsSCXFoch2S//3dTC8vWQuI+Kut7MAfc2+qd8rIFIvUWRX6DbvU17rTlspaUZGLL64
JcuoGg25HHIXzdEs3Xu0guUwPrD+/0NxG+vVvBLWAZhe1O7qYhEhS2vKnMxhyvsYboZaOd0Zmoba
X8z2aKkSES0MYGRMM7nKIZ1v7zBVyt/WtljzCyKjSUITR+8l8eqb3ubfqJsjxV0N5MIC9ERKiNAl
r/0bfosXrMwmbB2yIpXlCBkVe2N/EbHswARDL/2padx1KzRw16j8sijmFT8GyWyVVjMfHidTxIFo
P1CEc/QnzOLM/jdXm4rLfjbcYiSoRNxrS5MTXY/y1LRCVBGrKVup3D41/0nrQIO8iyNMiKWmrI2d
E+36GQ98SWTD09LxIReKDq8SkQKBKoSAiMp00ffV6s7+wWcazhRtxCnQAahboLef1guqo8a8+Vws
3S3J7WSzdmbf2/JYUrEzL/L2fz60NozuCKhEUISSWkSSC9OjgxbN4Vdrw/1mkZmhseZOl26G1ASp
8wgfwDH+J8Rpt/azOvo6KyM7P/bl1eRUKMOj0Y//z8TzHUUrEKZIuAtzF60GZY9GQj6axJjrsl8S
aUwaj53/5zAup8vO8gC+2OB3hp0aeKvktdBbVeYPlARt43yVNzFYUYJaagDYysfn5kiL3PbjyxMT
8kWi+P0vXh7BqJhr7WwFJKYp//xlGN1O8QTbNppJTugqu9EvUk4j+5ru+/OrOERsSIYB8+AvddyV
7yjC12xTSSV/mBK1i2dQp5pNBwtVW/hgz5r6jVqpDBBisA61iY618oW24RSq/H45DMwQHXt70kIu
qk+a9Pz7ZBOusn5ZMb/vCgZODCdbsoXriOjc4+J/+tcVx8a5WnB8gGo1d0FEpmNN96wpRhPZT3eV
WAdagIHyDNf1R6YVr1qezKoznyqBmyCVgLx+SXZ6tnQawrU/B9o1n1dR1KBFx/UKQY5Jc5+/ay7K
1F0ofqGsNlFgpQ6JrvEREVhYEQtpZjUDbu8hgd1Y7vsDWoxumkmjm/07fC7dgfxRvVqz7bT531qe
e2UZoIezsuVdkmeCraJYSztspmwrhOeBL46uS1kh2CHCG92JqsRJ3aFZ8rm6a5ZxZy22mzAbxUKs
REzF9S9wFxktIhSyD29iAi6lCryuR/xBpT4qcJ7xcCKsgiSMbW9QC7qtF/pIiQ7xnvdL+w9w/RiN
dNY1TiY3FDeSsVcQ4+koXoPPOAZsB/y8tz950bu1sMhgH1OQAwWLhdN11iELBr45rGPURp+0pmZB
CczhbWLd4Q+OszT2eNZhiWV7x8DP3wRMFFzSdTwlhgDEUfFVgq1oeVdwMTV03Vsu0b584Ft6rPN3
zXLErI9txnawJsH9NiEjNLLQEqaD2pKf1ifdyO/h5uhDqP80kP1EKU9k1h2h6H/MbgqD1g7VGqdq
5hRiGS1UqQlzUQ/xmZAJe+MKNY2HhdR0z/IjfL2q4DLixhBHBPt6fSasObD7uKV9z0sun9w8FreG
NWz0H+XYZumRM3g85Zc3MjMeNk9VUoODExF7I2PpJnRSh0V+jb7pDHFVtgUAOp+WVtRNh8bvLD7j
nNcqjAsMH6KO7gKMaPHs2PoXfwGz4odQcswWgqrHBQcQf2onb+nULWpdNfVWsGem8r2wvH4+nxhX
Uh2WojKcVf4JJAncmZpgmy6HiVsEMc+YT2Wp2Q+nbyZhmyai1rcCWCMJDw84tIQiKO7lpDyYFdO3
r0JYmFmxtLzmODrtTVHX4G/sqyG+/rvNRHVqO8YROxsUKBtNvcUBSEUJHFObGdj+BOb6gI957uqw
HDJXIkq+m7o2UpVsbWIENxagkbaYPA5TOd+i+eumEOvuBoPFxJ+iYgScOmfdaAeQYyeUolmkBQ+2
JYnK7/QMAqWytfNziGsKNCLQD4ERjBmJ97mWL7yBLys170IX3YdzTvkHgYJ4XPByW42F8YnyAnpN
c50nDoAB/e6LzoQ1Dq8UQpioQn4KrrQkmikRiDRZNO57sfDkxunINwa2WuJG1Vm0CpMUvsKtfnrU
gFotSRIh41TG0oY8lh9OtGbM1wS4I/b7wyG3mJzdL2br4ohp8chaDP2gQwE48aNj+dIQJhy2yNL0
cXLR4/nVpCULyo8A/UEYE8cZN/GReWqnHWt+zEqQsJ56JtZaPS8jGvI3sI8l9ey6zeQlyo7ULWoz
QWWzJYXweFEzlvZ767gvbJPgt2qV44NF+vPlAXRZiyO4WUlOy0y8ZcEgEs0q5fLJzumCekjjgmQX
cRrdYpfKWmuLjkXjCXAqIXFAYULVYQvtLIy709Q8CUnpoZEcuoI+SFIgE8NhpRyaijg7HNHox1gC
WQaDu7PSsV9wgbG0gesldGix3DJTbw7qQtVuNguwFeig0FPAQ9Xdortm2qy5U8KE8gNiPBkHwuIC
IJdccdNsDLtvYpefN7V3jQAujpqGQf91bUzc4SLT+xl8jOILNsZCx2QVctg7OVOoLRRWDIeWS6Vv
EH9De/r3EIL5IHf/CTbftSA2Gr8VP9k4jOh9OT7avXQ2VacRYS25R45giMbbKuONpCMWDjD3atxY
zHhIyzl6WJ3/p2OLM+biDiZXzSp8kWt3BznDJGEOYgpq0ZTPli9ETa7k7nRrI6JpB1hxvc7TC6YP
Axop17k1xe4HnIWo68lxPlX7UQsnK7pl9NriG7z/XGzG6qkhxJhmGg08vvws0ngd3QRsymaLDVqn
Rt0mlk4z7cQwpjRVLIn7coIsCWsJZz6l82iKALf45BJIvzlTsnPm8RTLAb3m2oMrxHBD1mVQlnih
3ctKHmv++OAoVtoxIgAHp7pZqZSo7hpUk1lgCNifyVs39d2t69N+0Ab5O630ymxiBwWKI1qNceii
fvfYu//6zMUeYKlgAZGSdqoohoNIbOZFJ3DLtNbZ/Hzr1JO49S6oaFURkkBVow8SvbTrS8fzItZy
3/w4Mahc7nn6yVSgik4NFLvZFDtOxRNyqk2BKoJAAQKPECkAVtaIjhxi1k+rn4NKaLU0cBoUPZRX
q7+Vn2WqIaU/ZZIq7hoodyqyEhnzRhbGXGps1GdPWwlgCF9ovjTWxxmkltDX34S6XyQthMX2Euj6
LgKWLAUoj3MUnpcxhMdAN6/nFY1Kw2AMd0EcM1dEa3zaNwibeLKAIOqevW50lKlqcfha+ajvSJqx
mOirq7nuWBkQxUFM46SnQR/+p1Ij32zjvRLXvuqMYWTGTDlDeDamU3TuYc/+i2njQD/YWDL1sWUY
qDAyy82ns4PotIDyJflDAwM+H8wO30D6EOMyAlNrNFO5rJuGse4AqoECdmuG8wVIahzfSLC9TA8u
eTVU0064hDmXHbi7ExjbjI1dHH92b5788t1tUYfwywEgnTWNTM6Ec7FnyAbG8jz/0JBAlfq9MgRl
U2KWcf411svYBAfgYnj4h/2FU8O1R61GNbzLeGGR2YS0rqof5qVPGW70efOTNYML0Gr1uGTVbqH0
jfbtrrtYrvX1NG2tIx/27VFZj+pPWM+WKKTFnN7KsLt9VhftCczJrXgs6PXWvM0H5BTB2K13rMHm
LnkqLt3mtXHqxbutCH0L+Pdyov3dwoJCfC35SHqpost0Ca4BeaT03nfuUH0YCFeVujED2KQwX3pB
RzNqjX2DqUCHUUdewBiVp8U5lStwIPvDRB3jaObM4T2Q4eHpWb5b7EO3Ef2IyE+0xBfCaoXbKM4p
Ysl+9sa/rzzlLHMuhb1MguZL43V9JExxUDZYp+Rh5cibA7RuokwBlEmfCL5ttRnEhv0oDhojF4cI
cnEHlJhrp6jWB+qgKW78Kpszg8KQ3urC/TolQduliTo8A0cMFLn3P1q8z45We3mirodADJ5YH7l2
QaEdBw85QmCPOSgV9NIImTb4qh0+RT7PICr4NUZf+0/R4C1/q5rJg4bSbN7Xko0beouIDQWeQlWr
bqMAlBRrhy7rmxyr54bTOeQHmLUJJmb3BeA1BITVPNzTsI8J9Wp1iwQWe2EhqhuO3q4vNBtDr9vr
U4jTbgAzAonTjyVE44lktQH4eE+247WvOId2yASX9asWx4oXzgwJyOVzsVqgWF33v+UDoy98EHhI
8xzn+K/qwQNE89Jn0xMS+ojanIl/WYtt4OJd8IKSho+bLOCJXP7i3f4DlPZpkPsMdNHl3IlWTF/H
rQtvbpFWNY/xnCPPsGEvfMr9fQRwg8zT4fuDypdx5tGHP1Ji1oMtxngO76a8j2hqcVcH+VddLQPj
xkDhYJZ7uyHPLKcZQQnxIyucriZTBllsiFz/XLylWBdO/VAgjahy6zFIcTYthcAAEIjI4rAPIL5w
ql+UVMij/USZ8Aqnl0Cd1YDs5gOSGPkUHcqECCDTV/lBHxnl01KIPGPLBiJ2CdDpOqF2btEvSYFM
hfTtGkWhZ9RUPqhh1pyWsIDjIP80AfPcNa4cdAq0cIIY+Fa1cf6934l5svaExPLMvaY2JcuUyT5c
DrYA8AVaJOPCFxcp4cvgusR2jAmMbK4GztTwGTh22UGBRlN8/fY8G7KhOXMp86zB/GD8F86/oKt4
L8LzqRvMRbQYm0d5lDOVj0pgEnw92xlqrQJLAFyE5G6BTqAsfdfBTj+ll2ksYyTUpCyIx3FoIpmZ
YzO+o+0FUfbY9c73mXj/6Bvl4QRDwKW1x1kD7MQzNrHX0uxzGafK5MzBcS93Cb5NyB9PFxSl+UhZ
QSBJa3w+M1j+UFQzjLiuRSeDVTjUf7x7Ff1mEwkZOx3AsLo5MXeuXEqGYiJvmronbA+d+0/IONwh
ANzyofpV8GHs1NItOotxZ8DY5ZdwoaSMeLkwVoSMQUNzZYB2M7g0vvPCqjNoY4jZsIeMhk+exFdy
MthVQPzkWNHcRHGzLc2aewQzI+k4CBtngEaOpaEy3DUol7Sew5MXavRknxioEuZkEhFQdRAxBjNW
rjV1KY2cwX1cF2N0GQaId6riQsz2SAj5a8NyIOShD1W+pKTUE9lr05ojBMWI2hEWYCJRdz076ruA
toTuRmKyQCS/D+W3YJeGUgsr3ahrQbT85cRZqvO6NW4v/sOFx5Y5OkgMLlb9SSLtqZnBwhgoiddZ
+1tfc9GPSOgxWE7HU0I9WR8GNfq0sR3iFtTmUluddU3PG/Bg3olrCzU/h3ItGunoD/Bmb4/+edB8
8Jz8P+NRaCOpOnPUt+SUh8pcJIhn/XwIdc4v86fnlKueg1qKCinXE4HLDFCtZYKYhNIcPQafcI2b
KspxyY4NFGyGYyTrzpY7FiIPWvxi6QFg8cfEXwfpdMttHbtv/4umII26pv7bYVwblN41ZQOCOTQY
V7TEMiNuW2tuhCuU4ynxXV2H+L+avbWzY/lQ3BOvAsPmvHjmWVOmkJpMsukVEKR9O9nCNzoduuwv
AUWd982Do3LHm15WjUpo4c/P5WOUiwjWCC9wyMxVrmS1TE17jRH8pC+YtfyqhhZr54cAz6mCEaLf
/ewjDYcW8AB4BAZ3+tRXLBBav5DYJGosQNVaBMNhUsReN7SWSjnfxNX5fXfFoBRGglOq0MrXh6gn
qSmB2I+6U2RxaCpWECSpdTa6WRMGSdA83VhN2F9nlYkQGNxWy4dkFaERpDgea6jnlZMD+D87Loy3
tLcNTwhvJkDHHdmwvw+lSppsH8ZMvNmA0Ji6FdplmpfM85o/8ReqBBNb9fKo1gm+i3XRwXTiQUWd
IDYRWZbkMV5cGRZdEEniI1ilVSib7dCi8kQhqyN0uR77c8k83D6tT+7AwVDs/Jz1Ph2kIAVPTJB8
1xGqdKliovBDWgb7mCKdY+/4CzBpFooBQx0J3KlpfmzBUhC3kXq2sZAA2vJz2m6f3WKowuFfz1rp
5nDO5iNrv+8Q3VLkxsy2JHJla0uCPOqedBVxIZvfZZzQ+6gh+vWUH/cNghyskBCIysyCyDLYIs9q
HJZ+Grv8+4HD7nPpCzZaL2LciWb0Zh8zSb/6Hc0DrNDR0cmo6Uy1iIps/gJNGZubnM8npu4tPCpK
Wra81146uZf/4jJqOSXpMzYLrg5B+G3P+eENm3z/kgC+Z5qWO4K0JDmc+T87TBlj95Ykc2x36MVp
uN10aheiTdyVEn7QfcCqlpQv0f5BQcVLXmUkbE0GIDe/08+7S4ri676gS1We9LF3Fprg1rZ6qWR0
jfyj/HJowJSY9EMyuF0OnhaoJLxTKdmwy/HJwVHyrmSVr+/iMg0dYnKaNftbKDFl06m0+NolJ72c
T8KZRAj6DTFy0s9jh4pIl4qy1Je36oHvZ0H3pLv2JQenlYDxxYyqxe+LE7DMf5a6lWhcleRyrZoU
Fw0D4ui3G6YXycodY55NGKkZYWGo9RnusoE5kMsbZslzJtSKqyMx2W21lKjGdV9Q5SkFV8+b4Kq0
Wz9/e5EmVMrfqjY/xUIlWxnmhxfZSkjuUVdrc1j+a3w4vw4ImSfO/BXQJSJdgA6rkjMwv9/FTaUh
nU51S8oP6GJ+iMa7RPkcjaZW1pU23KO1flAk70t+w8Gts17YliLNNVMp+dcfgZv31W2pCW1nj+al
wD27tRY1AN7hRzFd2uIHqtX8PkQaQQvnqM7jnWgXqlW2zB3mHVAJPqXCsBVlvWyjD05QM5kSSCGg
ueKnU3VySAbVjPXjshxuOPoeGbuwAfmpLq3gYIOu9ZjX+qB6DeHV7+7IaJ/aP39Ps4MZuBowZHp/
6zeMam2UXykAO0zYFCu85DET8KXfZH7HUvMoWMcmYluwPjp738/SoZrZQhmENuCVUdIT8CFnGEA4
4TE8a7Ok10AfxNT7VZ6Ppvwjraa9k4IAksuVokADsTxHNWsd90tz2xR7czBf/0g+fJGBmiU02zPd
my2iIiicsHsCON+XaKLoeoeD3KQucu1T69IDBmQ8U7KXJyfgyfQzFyd5ZA+GuyL3b15+S3vYSR4F
z0nSL8JDJZT3eCKUBjL85v9CPK+8cbYLhts19PkkaOrwz/4taiQSwgubJYKTFks4Vk7EYfkoQAjb
mV3CDofjS7zjQ6PBFj3QeP6DnAILUnng4/M+kupKSluEArROsQuctca+b1hEVlGOSdCgm4Wi9OGD
qupYbmd0+hCEGqJ9QEC/UYhtArRFNJpWjbYepJbJ5+47kqTXba2V523uPw0zF2bI8thbVa2rNh2D
B2QIxoVyhR9MclH2u8on2tPzg0cj/w4P5rfbl1vawvT4DxS8rYmmZcB0GRq1er3dXqpnVtS+iACr
LWDHJx74WRJ3q0ZGedKPYQzB7uHMTBvUh4VAOkr49rVt6g7Lo2nMD05zKpFN/wgSE3g+SCl+cu4z
6WKIWPGRSVBMNR/9MnFBgCasfeOnLnGlI6BRSnPMq177h0umQiMU7P87suUxpyRKGQr92Se6V1nn
1LcKE2A26x8/dL7pzl+qnT6ibaCr6kvnXW3L/uzm3ykOqV/mlXx46PqhLPttCaTXTzNyZo97VSPT
olKz1VBccKFhxO6DAnmOE/UfZ4xYvcvtb9LqmOtRpzAga9e12NIiej9UiMXE5udMp37YUrlfgqP9
grTjEcRtT9F1e4U+C2JY5ffQNue4GqRNgQex7yZoBJ8i05MaC7Ej7Mgj5DcGgIyGqCnoPvgnOPFh
Yn1mFYZ/nZGcuFJ6fzXmp2Zlo9Bg6r43G9LdFp1Wtn0i9+8M4F18jgkTXS3e3JaV6LQqMvtf0oPN
xel4RUF0HaRnwtO5W34VBwwkERVZRO8Npn3nlHjUSEg8e/aBmcLqx5966hfuYt3AFNxH/qKS3B3j
QDvqm2607VvfWZqRQiDpwLF8ev6Ds6VOzIYtHTZ9y+OpnDzWj5tJCaWvVWbft9cyniESo5uL3+4i
3ivTXiqkhCBRT2968x06m31u4a/5cqP2krFx9uW5Kjbo0nLZgDqOCKpbJBlmnfpXVLjItOkRJqmZ
S9oDdXlLQecZ+BlnFiPhr9B0IP58V8gJ4ThPmR46/MQGycuCBg4/rnyqU9x6grwyy62yDIfydhpB
ORppC2vXn4jIi+HbDXg8qvj7bXoP3TOfFEHUmvd8/Lv8yE+qhJf59ssQkPNUWYICJMkAn2BDYW9B
6bQ9/uaY3fWZodWN5/UFvaiNejvdUn2nLb7m+QWMZhHznbAXS5BycqMC/oC3A0KzvjCQabtNaFRp
Uk0lWljqRthkupwD0f3zuO8o/rUSX8wA7ZiODr7kMHr4uVBrcdz2eD2ZejN9I1KjQi9tqNNVxdD4
P7liarTOxvfL6p/FXzJIrDBzeXb2SIU9dsgGyKXjjZxPMBLqAzw3AEX619wV74B0y4btY+oUrETs
owCZ+H1iPYWnj55NPxhlFan6W5eP1Vyy7Bumq8Ol6GRW215qVKch9O4IIUAB0OteqwI6X2vJJt2Z
9AWE3hUKHQCoFYG8Y+RWqsjWUcIpY6YTBMmvHO8FB0R10RwpdYgkmSZw1k3dOvYyJn2AGydrQooh
cN8mUSf9oCdMFaaTGDFlzJErCFM1HH6Sx13jhs0hmNDRmBeG9KoX5LHUPlwBy9DJh2X1tjv8F03k
Ad5TjaoNxcqwQhJ9Y1oIgNuMuAlYuJfA6jFXDeWVxlfxRliMxo232sjfBwulPeAckWfUvQgD/Eiy
d+2nxK8gS3qeHrz6IN40uW1kK5E6ETEHwREJARyUs5yn3Fs89+awrusmURgWUoSnpQVKKqDIegD1
RO9PmS7sbFjGNiv9UPfRtR2B1MslodDmVn1EA3eGLDYK1RlxJPK3jOV5I3Q44JJOICXpj1BWAT9M
YJ98P6NJ2Rs8AAKzB2Z6rgM7/ZZDaZcnQ35+vVVRKc/vr2gCvD7QHqkzcLa2Ks2arpybUTsLzJl9
L0Y4krS9OcZeqgBHPTqVJr8IVIiw9kYwegmGglRb7xzqCOgMi0viTixU8YRK/rIekocpB5aupgQM
jVS2a8Xb9G5Ne+b8BSbw1+M9tFktAw+GRwq21ZPyNZWim9VnqoczOFyR3ldChYl9MKUcqB4YmGXa
beunxVZp7wj7zKSKydXIVgXDp29pPFBgYrguKhlfV10RnP6qEBdmRBo17zJsg6zeApwz9r2X6KfE
MNv7gzmMvlO6oOKTspGqgFMM6KtjpRZoT4J0U74c09pXE3SRVZfmxybnZ8UKFRB0bfPLf9Cxh0H8
H5SLkUZXUWLyjSv6Bmq/y8F5HGRWWWKe9lTkm9Tg8Mpd0ePTnHk4xCEfEIvIcC3gsh8QiL0wCw45
k1jcNv9HUSO6AKokwMyykvClovzQxnNYmsz8o9VzkR+fvsjrCwCmZIAOKdaNILUVyuMwe95H3LYS
BZDLU1UjpAJlhpZ5uWx6A7xqW1RBXduPR3F0S0ooEFgel+JD2UoB39uqXM686s4f4kGhDCv/QcR0
lM/kHX4Xn0Dcgipj57w5dY0HW3F4iEzNwIwrWHdqKrhuT/6NVvQSM1Q/5gZSnVYK3ATbM3AII4O5
AYxbb6BzrKJ2CS0CQoQ2woO39b0DNrkn/wPEqlALPt0dLf1IxtNeP4qYoJCj9lfjcXCvEXU04IkT
IRZOBn44p7iK/bd/vhtmKVQa4Gh3U6vx/lf035yu8NtIAUef4NjytSt+za+ff2cTXMczvLumwCq8
X+vi3fvJ90dygy/D/Nde5BDZ9nevlw4z+BXbLrMPMdT+S9E1Sya9mVa4O0IEIPh3gFB+7T3ZjTck
QpSTcFbmhFqE0XYcW2H82dNPaD1DHWJNL8mwWaH6tThWyLiFHxVyNthw/RIGoL1eCaTkUQcIAZQD
4qVh5Sm+JiGztC7Qxp4mqsG98lUy8H7OjiQTkR9aWg45nsK2ya2k2HgVmOqUtlTcvA2jGEioK+Fb
r8OxVg1dlOJr9v0kWFc85ZRmAjM2Vol9XJGFw0MHnox0qQXg5yJsn+A0Agbl9CDm0D3za/ZPSjAN
yhHvSCHCgD/AswdhSN5rv8wRVwpQbEH052mBW99hlp2bWBjhxgzuUEr4qGFbLS2Vi4gTqgBByRfo
n3TJ/m+p+OpNHVuhUYnAP1Q3raBCwq6howMnbTyAPuB5udwkJrUSdSv11qmNXwSfkjJPZmnCoT3W
Amxz4vPEIOe8iR/bYJ1w/Zy95SOSXHIqsXNDEgAvGjR62HnN5uQk3IqG+SvkkvwwIKdAj5CxpVcE
4hBDvglF9YWuywI7bSVC/5QHU4vX+sls215mhalIl8dGvV2EarpzDYmSjDf22WHGY+QFC0PRSM2x
nhb/Ow+Hfd1HKV3LxdyRQez56c/WU+/3s7F0AdxEpPl/dKUibdXOGhwtTM/7/mp/5ko4olY8U1P9
cnCpJSjXQwobemFmj/tUqHk2nmhZrePViIL2M6fp6/pF5vUWIDuVBwJ/6Px4OIsy5YN2TLFzg9Jt
LdHum1xFjHJtKs30SLmTBwOw0T1KbIkpJlak72qj5gbkDyEUB8tCwEVygGpeJQc4GZA2yqBYpJQd
unjE8JKb2AKedzlkKfm224WwgScXgLLuXFb9CuP2qclBFUviFhS5H90EYLpK1nfZ7rQh1UuuFlJ5
XzYNdlk+Od5DOzq9Ea9+XcrgQI7SDVDCjzE33ZGM5HcYG99naFkSlzHPxbq0gxS7Mpov4BgzimZf
on75Nlj6ioTwWeInSQFL0ZMgxmcRGzgv8TOydoX9cfG5LzpchfDE1zN6hhxhD+3yR6lL4eryZnTA
ZbNHbTB2tepc7AYRp9DbNjK+RG5g3gjqk3TmRjbHvhzvgYae4PLyLJP48N8siDQ33J9WAE/mZ8gQ
J1KfschcwX/Ov4WoBN0yTEfoBbHMZJ7aWc0S1tluy6bDF4agPJ4+SX6FrliVO7MLFa2lt7ySpLJw
Yp2ictqxNtppCgWS3fL0OegcDLuI+dBhXQRusIiQRMpllBV81S9Qri7ffaxzue7fM4I4fggYXJWX
kuCRlI1f4EgvSEY2kCmgPp/7LpZj4NR4duKLm/7M0de+Q2/aEM3rHc8uD9CDM1lw2tWSFEvK/ZpY
jCskF0GqXmuEEhsOnA6oCLs17Fym02bKsjgtvYn2D6pzzHdccK3AUUN7lKC+FuWk2iLxkDUE9g7V
HCUSgslJx1I6Yfaa21JB/D/atK3p2ulLlemVR+Dhkr5QtaCPj9e8vAD7EHPF0gYhIluaxTPDQ2UL
kNwQlvufyzjt1tWdhRR3neKfO3Y+Ee7hsjcgoJmBw7dOGD6h2kHjEyJckOixpOWdpfwfDxVL2YvC
GIxyYTxeqryccTLODXaiQ75+4ZrouFhguvc/yvTy5g37g+KATNDzIg6UzpO3o9LBGgsuydeGvS/G
uvtB/7pIgu2q9ydF1GoqcJ6dZ6Lu+3kV2tBNTt9BnWyKWrSmXulxmvCUDfxrVNqgn/zFWa90TKc0
nxphPoZ5Y9Q8BE4Pia2L/pyh/wZ8ysTX/0csdguoluw9OoM7oHWSMQFAofnN54YPI/JGX457mfMp
C7IeMI2WXPkTD93XtxWTfreelJgb8b156JJ0RfNO5ic4qAyZfs8Y+Y/j4Mw9brwRphkWVORIzoaN
mMUCQH8Ya6aM0+ZAzysfw1gfSeR1J/AKCTjzhqfFczqVBYw79ALtZ+IB1fiwvflA70SaKvFwlQLt
YwWAb0GzOcvTDnlfQzE0glb8M+l3HDg7rdasVvV1wmBUHlyHGkWE7LAExMBcdEr8ullC1+RdUBct
//h7WeJ8MBM8CWqXkrk8ofi+bpIMnpZH108DXihXHX9UfRixwRe7UG8c/qd4T0B5QkymkvJREcyc
Hbxvn3EehPp2AaUjkwLRYQp6PDqb1ge4mJqvKOH0EY54+TxAYAH11O8XQiZohI5ywPZNs35MF61k
mSUp/QROhgAZmHmdn15Q7VXmrLztcLMIjGFGg7jfr+vLxqkvRIkZQ5sAd88ImMO6Qr+H6yTsQBRQ
gIZGtghkPuRZzACQb8hzKIozOsuR8Dd5P9ik4FjEtToWr9nsEQUOnEdqIQT+M5Oo+uxS0Yz7nL1j
tXzWqG3lQkkN+/Xn/O1o3k5M0byxtVS4xkEVwVU1epJQ7y5PO2kc22wUCKoXkFwcgjM5kpulFGQx
1Y+MOKIvK1mvckg1DkEQngiqNqK1BzjUkPLGnc6M3DoYzZdFINq5Zh3cOrLQ5l37BVgkcPiA2gCC
NtnOyE3kuw0Gd0ZaAPLtJ8sYiNok6aSRHQySN51WXgl23QkBZVZJ2F6QDwZiiXZzUhCFeEHocwKq
R9ppLKRm334DcAzTTlBB3CgERMNR3s7gcNWoEhhAqZFWqYcT4pjZQeIuTwEq4tIp/obo3QTZCuGe
x4XGHO/uySUp7/J2xAg1fRwNT2ilbGLLX/nLa91jOd62ifuCzrhFxBmfVPzLXpNjV7qSR8MksvO9
T+fAv1X42eOlvNXmcZ2ngr4csKIAUGSQOS276URyJRK7uw/eRrcwluEcyHGTp2GUWOSZmJxc5Vyp
BWmYzin67d4NmnncV+bO443QsF0adz1Z4ZRShOEI6qsYuZsP0SIlS3VpaajKFasLajzYjGT89TMv
mTmohBb9N9tsrAQ6Sa8Jca3y0nBY5iAcd19byXkzJDOy+StkV/89C0zoh59MQ2rZwWtq/Ik3itp0
ctyFoslrnmIpWY3hkYPRC1PnsEoRTlBWOkazpQo+WiUrjMoltR8IRqPRz3W3RWkYVIHjJ0B5S56H
hG+6Jl6vpcYwK5iZbg4d9MCby0AOLKpbtCHfA58duS6fklFNwG2X4OVjCVVjAdAHJB5v9qI45WIA
61IVHyZqcrNneG6PbXEnKrOAf9g4xzzplvBZgHU4neQk3ISrmJC5Gi/lI4ATOq1n/FQlAfcNc6Tf
mRIaXhAN+K7qfIYBY30nN9lQVpFULwpxhJYzKPLSWtuEd99+Ht/ugqsbovkKTUK4eFRPkVzQTIeb
Y+8YIfw2hY/caW8sQrJtpAn8Oumuf2Lr+dswV9CRiFeQ0XMH9hDSgENk25rlQKasHYxj+e4haijl
qI9pOYXWzxaScU5IET6ujE2ULWlI7H4CRmu/igIOrZAGxIS80lOTi0mpio0a/E4Bx4Sp4eQot27+
+/qDhVJuJPPqnfVMvdVWIApifD2mR8iFOfLw7PWvNx83Snocu2yaghc/66mflBF/r1XFs5EKVM8N
2lUlE4uDn2uCakOttn9DbQF/ubyk5dpUd6qDxytiO0FZyaKCzj6b45aynHjrnWr5w+vDn2zmi11S
4Ox7iV2bIli4/zboWFjEKpfCA8rMII38MlefNfcXTDPKqUF7JwQsj2fIaGWi6iSmB0eOi3+QfGSe
x+BFc/2S+gIqfwkXt29LvSvdcszrMGLSJlNBa1x3UNzUXoZ5dV+gb4oMDs1mu/bpfoJWXKdewNOi
DYln/F2ZmAqraOB/ExBL7EM5+TSD9MsdQUBq1QDx/RgXfHL0qgZZ9vTpuQq2vmHGJ94IuFUkTfoU
D0OM8vZLsxD4NpiMBuB7+VBtM2nEo2HBh0YT9EHX5vT6SeP6KKUhCcxzeOCor53kjY+Igru0mGxb
IYPDf/q8gipB6iqNIred3sc/FtdnJHsmdg4LXVZ1L80po6zb+sbsNqcpYzGJHkmZybyXOuE4qMrH
pVWiQTCHhPCgxXVwvEJhBEvpDDupZvzP3I6eB021E5B9IAnuESjZpJ1BHwsCEfTfJTFk/myK10zi
TAznmvunfA3oNow0jVyLFeRQqjfx5CDjZyyPKPKz6TxupgyidcBZzdpxViKGK1nDCbbDtnfj6gwI
uHE7zslD1z/FbtjTUfjIg1miSRzDASshJjdUmEsdHZcP37gLGiSgBNa3mp/oGYETNhPgnv9h+c9T
J1AN9RMtF5MRJzJgSvHBXBR6rRAb+ZzVz7IICRpvSwL8khLovnptBnFNutehArwYuXQKg0FW2Qa3
OvxTE/XmbdkpnTqWKhF8wRDwV8YB3KILxZUqi5rsXSr6LsF50gMLPjFHSH1sK6acqBCIT/1cjJou
R3FYrUFHSdC7XzgwqSg44L3R35m8Jhyk2PLZYCOl6vty/bF10tcVGMmGwczoQGNJAoxJWjxi0/f8
pDsDZ1c+yv0a1DhQPhC0yN+MVTqwzyLDO1BcN5Yn6B7g33jhCteVCd4hMr5zAhj1QhVMWMV/qjTZ
jzh3LxF5M8uQxROg+5LK2qYkFtGIAxYwRDcXAk1iGVuQadBvLPsu+Ye33XDC20JkffDCbrwwvQ0W
MHEzmaUfDLbdV4ggybn3NkfYh7dGpfRGX4CMCC98WBTlRVdhnoExhy68rvWisewtvcFxJtMbhMjq
fdSebkdKOJepQ0ZXMqaDxWcnYrfuTrUYXnAQCN/eBC1KbGE29t4zSahunE2ce+cXM9FK9thlBM2u
TFkmpY2YuzYKEjuXzs9yIU3xHtSwwRqkZ5Vx1IHTdIusHJ0OagfYKpTE3/EhWp/lBn5XMPYhVY4x
Qqfy5R5JrprMSgK+QPZBMK0iSQlEA79vKuGoTQ6T6cEP3AC363XG6/K8hQ4lAezj9qiSCtHcXvTU
zL/+xdUZaTjxd6QIYHjX7y6N/eNZy48zgS8fUOoS5zz9EzSgicrHDqwBVgHZQVdIf201+mJs5X2S
gXmezX6BBaCgO7cu34Ctn2/tMj6fxjbOUUTw8YobAzLtuW+o+zHHodnL1FWPmdkk9rKQe7c3U9Io
m86tGcaTkoHSvjBuV3yKiVmEeciMx4J13P3VX+vP3JVPJFGwqlsr/AKQZl6o35uSLMtDe7gdfCAY
l+q/Alw9gw2g67JHrKuYr2YHBu8g9iZxuOkn3kMpO0pzMf8iLJqR45GjA8KCJEiumRcpGkY2ZU2O
0wmYflYHYLMycGoWzmwdWg63urnjti28e1Df3Of5ohMTj7eN3UyNBZ2BnL00uGHOvx2mgn1anjBq
ZL5uLP/X92/BLCwGfSVYQRrjdXIDP74yaJVE6+KrTWCRFLP1/Ew/7AdrAyvuWGTooXvuDrYCCaFj
5HrQHQ3baYwv8psMmQs4gx+YAB2xzPu4+/gogAES7W89OY1ydhlBL1q21NR6C411L+i552jmf24e
7zqN+vYcUvIjvZEoAczJU+w0DUj/Cb+GpFkpGmwlEv0ZiMolR68IZLBPHt3dtQL4yIMEQzka0Xx9
S4PrvoIzODxL9Dt/lgBrAWFLEIfr1K+Xpe2q8yqTSbAe3KnePgf2OeVG728A285Y4TyAuzOrlx1S
FHqbH6iFvb/65b8tbiI8Nz2VTUh5pEGmJoclDT5MiR7XZy/cWsE/00+ovmI6vJcszGEhOVxBb9d3
ygudNtZK4CemA6Fl6ewlW/tT7oBeim1+16ZNb4q5TdqbWnf1hPIhhQ9vXX8NShuyUtMBXlJZY6y/
aVNBG7XCkm9sV9dd3/vagXOq5rzHjDLFqHFDBOrUFq+DCro6iwM1VA4lTmHg8UkvbK7SWq8F6yLG
7PYjavwmG1lU7Axfpu+/XStHHSdbefWlK3HEWCSWC6yWhFMJ9ZcI9Nb+AqcPoYTZ80oXfhsn6PWH
9+Z7kcmEHGR6KbA10o4vUQZKlYTuLG4UmkCd5M3YKANG7Jpu11yUWs7wWTP+3iQF6InfL8qr4w/d
jx0ID9Q8vzRQINSsji5qqmwm3qIl6Yd528W8I9GmiqW5YsrcBYo5tNB5tmexV1ieUhLcuVCjzU/s
9P5ShD8JzZ0PbY7V1fztaVkQLUPiZ+zcN0NDcW8b/dtsiV+Ev7vCrWqTiAZ26ursWqT5PC4XCYk+
rBzqSusoDYwIqRQYnrH4R/HELvCSn9uPXelI4CDSHSUPZYouRepPvcWbjzjSfiCoimZius+WeIxo
/VnJ8pQCKz+2t9k3u7r/wQGhIBTXSUAAxhAiQs6/O1uTmLgXEXrRTFmWszatn7TpaWoQKe+7Xps3
A/Tl2gPbmXEE92dKWJtWIEC5E9ctc2r++iEYIUYOLTzQN1zEEhjyUhdkHI8SkU7RH1eUxYtwSqRu
RBvHYNVtXcflpfV1vvzCmVO4i1mArKtca8Aatjqbn5xoZiDfhkyEPBZVK/FcXEr5TDpG8BpYgZZt
d/V1SJ7foyCnr6EdIzXdOWkqAJbfuQr3z7BykFC90Fqe3W1C40Nl3D3d3LL5sdJUbctjWZRPYKHV
6LnJIwxem+XKDTXQqsOXIeYr3lh6czUxDVVKpbKtmFDtoKJCToD57D2bLlkbmw9pHEoOr3iYhLWi
wnvvOiPSuT2oEkcLHqnm4vFwj4M3r8kPmeoXFYS2LPFSd6BC+BYkwCFRiWotQxM5doU+VPTwMr6N
/JMsqqwO0UxOO8Q/EouU8haW26y6+zPljjtq2tVPnBZsH5VPkk+XUWD2zkgfKtfvfnBUvwkK/3cJ
XDwhgVL5od7cwFAdyWjThqzFjfwvubAmBw9BB3a8ZuZa2qxTHW1qksRiNZ7jimFgz+e56lBupjGj
5VE9Ro/vbyXVG7Pzw1KwMc5CSysWdzPmr/MWMSy7P9CKLWEUfdJDQoeR8l33ijXpmt0GjKup95Xc
F4rVz/xbrDofk7XcmYr8h0Hm9p+Za9YLw/IWUD9jQ/lnH57qMU4yEdQ3lLca+9Jo88PCaLNccjqG
OP8MlYbveag1W5Ctqjh7JbXFolGH4yiLieqewMukSHFfSs01+MIe4aKkYru3dM1ouHXCJS4YLDC6
e0ptVv6UBi8uFI3R8ukkbd7lT1Z+pBPfuoyxWvTo0oJXAiC79E+50ESKyVR4aMEN1HEEIJkcYKpM
Y2CH59EPibdHhnu4MGEQDgWvKyQvzc35FiNYHq/xawF87uxFa90DSuTO20Y9OofPjseoAsJmA17p
QEHoYe9SUP+CWs2wggnoaOThzOkM5NmbScQG7ASjoeNdm5C3HWVT959AJ7eCkUieRaQmBA1yJwFN
oOw6nXIZbR+tNaFQmkmPlfJyXVugKpMjTJAiMpXv3Pg7Vj1w0afVgBOj7+FwGu8RKhuihaDB/9BI
12i8r2pHXbwKzL35dIXq1MUq3BmI6VLPro1tf+JpGCyPzPE2LiQAmEF7QiaA7+MRUcaOpWGW5laO
s/jgG1HWl/oTUU42tunX8/YMssdQFOzbOrYrvjRrEayD3lUewUDei6j6LbfSAffciwkv75FfD/7U
ORy9Mwq18eB2VAFhClmXv6C0dggvcxIdT1ky8k5T/x/nNB61NTOYW4QLVkcljgrzfnP42AphxSmv
q2ju2qL4eGu3PKqLCBR/3AaamKeyP97BuBWFWW4WWmu0nRwY/iF0GIMt+54gPtsRovs2/5w8NTXd
MW1jspYCc2mY0BkoFLndD3wODcBCmsVuDtX5bOpQGPp4n2CW1RWqWrwmGM+6ojvlFOzwaeMWXhGY
KAfvwDfZiaAgqKk9bVtrQLrCVObAhV/ndARmTp9ryQ3t2rNl7cbs8lmZ0oCOby2xjPc/qVE7jmlN
4EmuGrQpJokRmyPK6kSk5kmlQVB7j5Zr6U2E+AOiZVNqoLJlM2imM//PEqidkdz9pAexJN9Y5OBC
4rXwieXk8ue5ccscwHILKQkxDWDz88l0opB6625FzLEqvF7EQe2WIw94xk4NOXPhODOP7vus1QXX
wugNQVLPMGEhy+Sjb5S5cRPntr0Uvq6wg3jMIbjilA5bJgiMcZZx1ifHyP9C/hzNcFskz7QDqm9C
UedPAZGM5uJnvaOkEjONNmjhIzOZjVA+DqFbFUL2C+y1YNQqRzXqPwmIPq27Dk97az4bsTLubEqJ
HtpqfP+MNjgdrPaEpHQ3F8adIQtQXrE50n0FfR9qcUJosVi9xWd99pUkT8AXr2wRIZuAEcT1E+yh
Jas7/zG2kDl8PMHqtLhWhfEx1xiemgGW7bCaKmW2nq3bpAMRrmlnEeA/HkAAt0amESPgeS1ELgUw
CpY/Fu7ErxZqsV70UaRkq6NI/G/3OOHSo9ICpzRsIq0/0lYzF0/4052lItPBC3C/fWBRWfmuzKsV
DGGc8+GTJZFQvA+kOcFYNu/4Dk0DpLP/laZONn0vXd/iIBbYuUL7hXeXUJ/iVq5KSRBnDzgvEzko
RTAftkDNaiBRsHGaCon81pGpdcvEQYTjIrsyJ4BlA6QcIXmlwjjQq8jyg0reaax0ObVGQeTbf3fR
saogpHKFa50H3c5Z7dJmCl11r8FtmOLVghDvXzqiAU+oeOvnrCKPLaaL5I40A793cIb/p7KiceRU
43fMjn3mxfR+EJ59NNVPQ1sCUrS/SB9vdfr1tjZkArjtMt0oewlTShV/QYerwLtXwAnjbgx0kDSv
Pjb5u1usZAgnS3wa7tKtP4yc4xnWz8jFrEV0E9uZG8Btf3gTIsU03U/W3TVsvD4KqDKfvg+sNYEn
PFoQJcJAZo4odTA4V4eJkAU3dboiGccrmZ6qC6tn5o9v/uLocoYErftNKytnPD31EDVrfIM/R6AX
DpIJuJfKKl/yYg5RMsRBCpUNloP3CT6oiC2yseIxaqkIibXWrtzcGRNWOIP4M44C4VYuD2VKGo7S
LeVR2Xead3VxLuE9drvIqPpr9tSYOx2hMDyTPee0kL3pCs6h3vCnH9Et3p/83Yc6u2+hBAZT4JOL
1ck2m3fjQbf6pyay+hSPSc+tZGsdr/x1/k4WSCz6B1wyOQw9BtpYrdU+Tl8Lh69nHwuO05PrFr46
HQ9ThtSvv1vVm+eRK16EYRKKFJY7d0JWWL/X2flwT1bYyCKMbjZFTfWas2btOy1ZRB8GlmWGSlMT
pUOsKLwyUcFH/YgD1nyUx+XkNQo99Wotzpoa/r0zQndCB+mdopSCdk5OBd62mJZo5kNTGTRJ/W61
foLgv99+nUyw7JUQAQxFqvuLyUg3tEBM0KW/Yn1BsBYhVi0Vs+E8+aivJv2pzkurTtrg/NC6sC9F
Y+MyvKGsGtNXgowbDuFBP3uLwDiO0Q18bCjiNMvukO6HoataN6hjZf+udFHZFaDgkLgx5BaaK3FQ
pwpngEn6oSqd52pkW+i2nVLnG4YzEsHEeo/eIQggElbcZVzBgbHW3M9lHgHV/MLbtXFkNjQ4HpqV
JftF1UginjMACMCf7bRxiPS5rw2S1Li0B/dVgXNckzToS6wL/UEH/N4jA6RSnKdbPxYYZig7YO5I
5w0C+KNm/MSDrH0KasIR8XQ3quaBcuV8ZFVrCfNCGWbqgnQwekq5G4NEWTQAbb33gy/bZpbnAsaU
HMznBGgvKfuCtg6R45wI29TC/XUh3qX0mjbGHjG4DZbaetz4AAh1pbR8ugfGnnA6wbmq6yPHQR3E
CRCuMyP8nsphbN6W5gDy98RyNhSMIpjvW0F+xbv1Kpl7r0kScGMRR67nefarvVRHe7LZEThAAFCU
j9sBDfBl/jBFB54a3L8MOf3gVCTGRJKt25i6YGp4pdH7FqjjUCMM7LrGMsGjEXwJQ32rzLinVoGG
F77YhKnNl9tmbZRJJnnENGEWi297kd99mutZMLZArpoLArMcJTORbEGzDNf6FfSX4iGVvVRK+SeQ
TYefBNp8SZF3usqtcNLna+SwTcLqzSuCp9AMUS4zLhTZE2bxLfLQ7BHZgtxaIu9vuo3SvFhotivO
Ntjz1M2EE1lBeWDAaMaRLhT+RWQLTBVCYVNheAsY6ls6bUTPBskVsxQJ4KeCy3tHKjawqNVDPvlC
8OtLtAp3SAUyQYpubOUu5LngWvaHsJ+yGvch94XjT6I4VMQrHFHfTWSTP1wvTLgk7adQEgJb3Ttl
lDS7avR6HEGRE0c5SdMEk5Tdp6X+qw1XEIvnapLuBQ86rtgcIk26BVuNBCFmPgqMLzciXps/RXvi
/UPt/69sxup+aFDnnYVvQquNlIhlt1pbFQfRG61GndBe/eY+a/IY4kNUADDilWXmTBF1XAvFyJU8
jyTwrcPw108OQzO/G3SALH/pTe63Eh4mAI5R8XJIeGjPlNXF9GRQcxaiPWWD2LRuWJKUvgStLGtr
/Chu1dGxlN3/Uoha98RIgdtrd1SZrixSkkt1/2a9aJBTw4Gy8VQLpmy7o3ClDaeQ0X3hL9lEv3gC
qpp4uckwF5GkxOPfsxSMBinXeoUfvMN7BxRXknv1+7UaYsrZs/t261fp4q88gNHdB5XXPwcf8Grk
z0q+Ss5aq4evZNJEeeXMY309xmUP6j3gncK8z3qFiXZm2zZ8+WnZ3e4xhVysfcYGWGNBbAKy0/P5
V1qGodajfZG/9ERUqZTwJfehRVK99gZdMnhvnFRpi/+SOCTjQGAqIeqQDXAdKDmb4Vc0obotQ25l
OlVrbzkL3BdgO8d+PtFyWzE9V16p76u4EychezZ2a8VP2rDgNsAgqa3lFx0XTG5nieL/oe85kNbu
+aCUMgYwvjvJo837RHnQg40Dj/AJp6T1IV8wpv26U4v5ZKHAzYvqjX6negIJiXiZzf0RasTX6UkD
qlSGrpj9zy2d7ZV5o97x/XzbpBPFRRIFXkDkG4pdAkj7SQeuz9P4gDyIalijPBxz/DVHcUMguXMH
vx3+VSCppzKjrgD8arqgKslnqHjHEMvYHZSQG20Wfg+wJmNo0THLHKchuPFZrKYiiXighobIM//s
GD3kpWX8oOlAVPIlNyx35h8sUOgWqSEyMA5yZREX1mRRFzs0Fwy1o05zJ+MsPKakRMBmWsndpvx2
PqSxfDJgDiEt5AqR8Wh+Zs0WBaHPanJZsKUQ1lS/te4xY3e/y3BizIhOlaKYhzdmuKHpzUVCD8VE
2TFJOqbwMZ1TJhtcWQQ/zi6Feignak7kCirTqI+HuXwc1fHULkd0witCGe9ybwznYwXdgz+7BhFw
xbuB6jToHcYB8qhGh+iiBd/ODRQf2DjC6QpCI6Rg8sAa9Y7/M4Bvw66ENUXarlN5X3Mye8Nne1TK
FudRgFHUnYrdv4e8MctWvLYXzRWW2amIe6k2N/s3wLyla4YdEMzabfg7NSmXT1P5rNhWCP0V33QO
HcCebhXcL6Iu19eZoeO0w22Lyor/f+MjQ2jmLzT1SkgALW3mlXDowXQyoek1oXGreDWwkrewOnP2
8DelgWJoQ+vdMn/xzOYOAku4XJ+ISyZpibPUBiX/3AiM+1fuNHc0wvmDDGQPjog9jKgMY7zLCVO1
9TsuW+2BYeKab9mx09+0NunEEyoTAc4m1Jk64p+6hMpNu+19lBENzBiaeGiEAnB6w5m5xVCIXLL/
4vkvsdlfYnwCht3X50bbTDkxv17TfmT8tK7nikANCBmcsto37Psfqt8N4awlpPKcLTqfmwFvU8mb
Rvz3Sgm+C1ckN0KLP5K8w59eZ2VMF0Wf3pkUAWzwl1ezTU9ZN0Uop5Vdi2TDPdr9HWOJm4bjOxz8
dCPFUBlV0PmQvzhjBdSk8zwnizY7n208BzbjnnZ1Wsd+PYVqWIPeKyAcykBeqTL/TyC6z+823Cl0
/jVolHdiG/0YBVddw0WV40pznvd+j0DKWlmhFd71GUWndEJDOUufmMfQSzeldmGic3qOzFIDMhiP
oyLPYqVP8Q/iXD9ME8lf9N5bnDBL4CK1lHDhbr80BoMJs6itl4ofGYt9Cd50IubywvtCNHrude8s
OZTHMWnEjWHcrQvEo+OC/nWHx7nNeORSne5HPImvY1wEBMVc92mCt7A12F+NvpjUlOYCtfWRfKip
euonftWETjInEJ9hTKBZFIPdimVg5SBI04FobDGVDVJ1KpeLyCCQuRFwDepCHPILrrmCfLs5cjUv
LtjhiwFLF/pQEHh/I1VCmHe12wA/LI9Av3GerWb5txUbL6yqM7USHPLNpycODIf3H/YE9ksXgayB
WS/bSzPJGBrvlaWzDxaVE2wxrD6zr+Vv395gtTyZ47VxINz0M119w0CFqRR2XaTzYsQg1JQw69xE
Vp5tAArMSVSxXfJsyuCd7GcJkkfogFrdRPpZJA7duIhBxwD665klR2UHo5hqiWtDbMiuuxKaxmiF
zZL2ZAhkXchFaLOV3/JBfRZSC8X9mttadgeTbnUOJIe187L9fssMGGzvbSWDGcg9Gbky+j9GQ6N1
264CRYZtx/HU0wAXMdjsxATHI4N/UEXBsgLkqfqPqLMaDiRwiXNrjgOy2d9EL9dVJAeIE1pjzPXT
XdCgYyMps2AFnmLOTBkNzppjY7ksukIRGjWmWQuHwWZdeWOJCgTIxYdDe1nJnxgFIZLWT+x+Ycqy
MEpYaJSa8/WPPyTWG4rUx+Qdwt5Pgizy68GgZ+t4ZnSjTwej6qe6v3eQ97fmDqsLfKdVZ4g7inWO
GaOcU87zDBoxtGB4r8GhQeYdICyXW7/t9hxxi/uNg7xVqfZ+W/jLPres7OVzkk9nzcoUkcmAK4j+
MOeVSFrsRBbjr5mDdYkjEdiV9TVEytPC+MyuTTcgPxBCFIPhZIM9tX84lOC+dFA6IGZenPmb8Xsn
mz6dbkLq9ZK9IMstiVaqA2X/B6MC+SUIU1+Y8axOjgFpP+ljLtdB495+f3FqMRWvnti+Hp3bDh3Q
SAE+VJ/eMSGTukS2qtBm6zNEGIoCsjtb49cnHm2QxULZrbyjJW7GVhdYiE6OBk83hStwuCh3kaNG
gpwD9O/wWUvPDPG/vFt36a1+GbTU9O6VfuPuGjNoujIMcGdQL5NWOGhiA36RKRyO4/TBcJEGV9gq
oRcS22gCFAeqhxk7a611tRXUCFyoruriyEM+wQZRQvieoMGiKP6gciAPCBo0H/yVsevyjsy2/MKn
oTkKj90docOdeuDN52Z2L2fKkei1RYpfUs3VsddHS4I1lXMP9zKwrlizCp0Z8qgY9BtQAuSo1ERq
G5LMmt9qykU/wN33dzbrIL3ngurF474OO4EtJ6+iC6pN2vy8x7cKkM7x5iSrs8ukDtbJwoemvCIB
5+5hZQ1bZETA6DJxtcmQCUzhLvgaDT54NEKfdBdJKbkMYJEiiIaAbt0FqUtGt3j9cSUytEi3LkXI
Ff6E3fPxMV7u5v3UKauov8/V3MAkIBiKTYOTwGe710rg8UXDzDJFJOn0ojtw+Vgin2SLo/0eoLCA
vgTjRAT1eM8B6th3tpN8D34jgqL1dItTz6a0wYug6RA8aUxRKXbxQKpCd3tz6lKe4aDWC8ldvkFz
8H6Q6uvgyi6sXzGBLWyv0JHrfwYiV7rOLX134wFtTVm245u5Q87yYj5szp+grdVX+LILMrZbib/y
uvSAvpEqFWvvlKngHAatkx+RZI1xKBH8Y/Y/vZBgUaxbVs0Ui9+P3256mRyDQvUtj5R4Ajff2yDF
eV4TrcydGFfcLUET0YXsokG6byl34GESMwMkx28W/Lg5k0//4eKfAMLjo4bR+wBcKskDk92szn96
UprOBcc878mVyOthagvWRDUUgcr2onQD2GjUA/CMCD5yNquSeHF/4uIp+ERHf8+jF4xw8YMdT/sj
k/Xzjq29dFJvchvOhpXrLj49kBdcoNacejfyFmBYzlxXTZ/G2i6lmc0kW4S8Rs3Ukk6mME0GTchs
AhuwDkiRDcEbgkU5DbAdYEDrdszPTIpIO9I7+VIEUK6fylnkHXVq5ea1mI7uf1US/SIQeNY3TohI
Sx3nA0jgvBvJ1L0fYV8K/uE/sc+h/RtiUEfqtKFNSJyo2srp7sHgmOyEI/spBe6aq1bU51w/+QBI
mfY70+cjOa8P/okqmPRPS8c/GUHFBZn2NWklqQwMkTb1LR88KkKdTi4jzMHGbruVuphXckzNCtCp
DBT8BHihkxWXD84daznK0yvRTF/tBW3btT8ftVgoBGj3kL1Th4GgWspE+EcH7zNWX5mnXyR5byPO
oj408hmBl7Hzi7Mkkf8q2gTtTAMyqUNup2krg+IqVVSsfMH7H6ITiudftDPBwa9jQEcTgkEiAJEh
52jTQHHUSFIhMkLCEnGCLDB2h4vHjCwllUnhXUPhrrHLUk8YC/XkdiTxOy4W3if3sUzyjO2CAP8o
I9FJFb+oTdlq5J1OH7aRC/ugy2R10725DVoIWRicydHJz5AbDtY7a/TBIs2GoCoJ+jlY11s6PJZi
3OLEqTrXwyqAV3VfFi8L6d6sJn5rvVcGvFCl5Vy9M8BIZv33qz6F27EZJMVWvxtTcoOuxjONil4z
1KJ4AKZ63+oiL3h3Wbp73C9QvKvtsRfkccXmb5uy/mw25jIuXxDChAAOLZ7osqb25hs7dEa9+mWD
Ke+lcqAICmE/7hDnkwpIqUkEkP7DOoWD7WW5qbZzLxDGet9skV/XwTLKQz+7871kes5Hj5UJ+MqO
j3K1WWYjOwEVOsmWtRlgNChPBFPMvZgDCyuwa5ecLjIQlEuKbQPMcH3au34cArrI7bHgdq/OJLuO
oePQ8I7B4I5GatkP4tg0LCx/kC7YYXndKU+mKFVug6MmLKBx2uqapD7wiY5AUM6ft+B7xibmmwdU
EtAWqCphMYUp2MH3JrpfEKNMp/vEczVAv3BTZK87r4jsPIOt5PjDs7tMnJ1tW1QSwfPp1esOWjLs
xY4i7pa9JjEG4bsG30/PY1ryWQXXPR6rGv3FRimhPljBzzR68tNpfRaC/9m75fhrU/OK648NKI3l
bGmvTmbO5IA1YSqNcOy59BTOdlYEinqeIMBNU1MdzQnUDd89vjsNE5LFMyjWTXoswsVjQgsqGQSf
kKS2ficaHU5SKBU0XvCQ6i4P4zY/JH2+aajfdouXYUUZmMZz25x+/a9IK4Q/OyV7TpG3YYzLg5PB
sMLGMcuNjUeiUr36nQwFyl12jwtO4QeokdJY9sUOLJF0K6vALwcxQLgcbw0bDKPoDUPNBdlaVafO
9xq6qE7Yt6sYvJIA++8As7aOXzI3peOhnlhIQ2Rm/kEe2i3nZ20focqhvihDqEfsgwQiItrJeZpF
QIqhX+nNtwV6SGzzuulkC7qRNn54zgnZUGdbbCl+zPBLQevQAUfpqtp+oDi4WJfjmGbT45xEttE/
x+r4yenNgWN4EMpYEe+9xCmeJF7LX2ZAY8C4oOS4DMtMJNPHOvhOI9PhcTm3Hp6rMz3mmnVvMh1Z
BOhnHKuGn95/Dyq8gsjjSFe+zkYaB9x+D+aTSbazi/2wvGYhs66EHquJtX5lTLL7gCf973pMs+V3
I95pyAoxys6BNYkrXODs2SXNABHLt+24ihiSuqe34DhZNPgXP+fbgMGZbARtAGIbkZfojzHe6B9H
LP+/Vh+RqPKCGF9cTaKdLvkd5zqkZ0cq7EqIDRPf/Y0Lnv2TZImu9F1s/6jelVTSWBQxyqMriS5X
RdenRwzohXpHp+uS2tU1J0bF0ec0jRtsPhbnEGXsp8R2nggehX76pnK6E+nknXa2yiIAUzs+GIg+
2Hb2pKfenJyhP/Sz+kjIMX51fDFuQN/1kgmDa8326kJGAd5S2kBqHC0gpVDBNLhHbcncEHeWUm9+
LNpbhuWHPfQXv7pYnPj4CszPfSHIvb9zGGhViEWtZ1O1QW03m6t+pB6ee+6BGdqHfwD9mJEaLeBl
HAyP/NexPDvzO6tJlHcUqV1CEkDIrpW4yoV2J7bSlC5qVsrbjspSjwJauL8GV8w7VxETgZG44xaQ
X1WweQnsKKSt1BnFqxB0FzaytfEzdY/BodRupIJhtSM85f5mW5iqrt1p3l7n7bVPwRnKHTRxGt/c
RakpqbId1574lUZm+Z63EBVztAmHFG8Ge5lP8Z7R2an8GWoGYD8FGm4Z3ec1a/P3/+NZ1LWq+9aZ
RLSrEAksIAsxEt9V2MiT3OtjyHg7w/u/qp/7cLmM9QJDFJG+/NHQSbMDlb+zlfamOuvFA6OmtU8Y
ndSvcgTmyEuKNjb703vVeEChAjzhiAoCiHsen5BYa04zE+9WgBjERy9BW27+kJqhncmEPTf+G0Nf
gMea2jFr8ZckbDiWG+9mQHdFilNbuOPFewMxSvDURZmv2eYK1qMInOJCQBniDFLy809A8L7BUmE8
wsc5bhP97nmWKRwDCW42GQwgduHO49kLpcp6HL2zIrw6uKQG3LOWc1c1awF9uPbcDEePH3Y0YQvW
jcK3I9q0Ddl01Euse72oOyVP3qVc6Kl2XY/ufjFT8xlk3xKp3ysabhTUO9TokQnu63gjNvbijg3a
68b2XM7wd2lt6r9ukvGKrUl5uRd2fhl70dzTESwGNhbfBXLo0boEkwfTpX786U3gZSpPgLSHQ0Is
yeFej1dv3RRoAQjJXeTLIqBnaKm9q9942MoIFFD2Uw/mSN1a21r9VTPPwiq6WbIz9b9mp5EqOKcv
YgGpTx0vl6JNbq+KRwGs6ACJyIuGvx7z4lXCft2lhI6npYePSjsWC3zvL35zb504zM8J3FbFRnXF
GBfhcl8D+nQHvTm1I7IxFJCyR6VDTjoM56up1VVkEG0i7c6sBuT4hZHrT6W9vMlrUCI19C5kfWGR
BBhFNL5fhXVV/aIplT9CYFWxmD0esg7qmQ8kQx0D2pFESqOPJgP+z1lJZatF17QBfDO1dhvwVdYl
FQNYgU5gXBBK71zSNCSoYNLj9U4G+Y1GT5GB7T5uAqhx4L6O2Z9flDy+C8aqOe46Dtf6pnDW7dCi
5ZSFWc7smbzCfHpnR2cblEjhiT+nDxyaPDdTQohUqFOSkOsjE/e3X9nSTs/aoXIxG0Mt4JSuwFBo
y74uYdgY6g9HifF907LTIvdPEGrr4rvn+TnFgPLOT9Wxb5/hu8bw4mZyZ8hn+8SuEddChBguqpel
LKf4sL89nDVvejoCPERyIaIu23y2NateIqH4umykEhEvY+1zkm4e0CwCdcFmCx6vP3LFxGq3tcaM
79jY0Cp1ZN/r+zrNKLZiznYlK2AQ3rko/ud87KKsgjrgHtBqxYW1Q+Ds++BZ6R7pvZZWU3Djr3TI
VjVFwTHaYbre7jHGP1Tgu761uGEsMLyxwa5dOiKWvBpOcDJzj+/d4nE/8+3u6X5O4ZMPpxdp1S1A
+nAHr/ysC2tVhZ23Aaz54gAicGKoooETWNmkuUl4xAIgMZREzshV8xNAnjA7rCI/p5WgjqdHyS19
oNtA9qFzB6SfDJzNlH0Wic/gUJmaTSE7aVTvc9cBcMMZnqskewRWCMe60MiMqpSrEn6wkM+9HsRs
8jeia86i3Kq0rKuJucMrFVwAfLyQ4ymWsV0xr1zSGmSMRV6AUzB6NYg9Ux6iJxZLhfxw5zZyYfgq
mc00sFO+wMw2Pl2rIixCpfJ8dI38nv2PVs6zUimHFPg1KdqWHfaQtAPrn1AIwAEy7DJSUh0s8jIg
TlHA1eaWYfMztQTlqoPGXSgxq3udY0KO7PBaqqouDdR3sUo7VvLYTp7lOuRHOS66tIHM0TbMcluu
eZu/Z2esZl0X6O+SNaMMq3jzdOKmlpwcsoPQ5EXUIEY0H7ROo0HCcqutlsVr8LGIqJMTS4qdbjyQ
pIwyPBDVgNiJTm8DCe59iNgEl5t01CtwrA4yxFlC4Ai93JWQ4YC3bVHfy4FFQZjKpQyeuJXIgI1J
3XLeO9v3bhFIffYxJd0gdcX53SsIptQ14sBfoNPen4jJbyC/0DBU/ck5c5qmeg652+wkPcrJD1kY
wR8W8O+CuX/1YAVGF6tGPHg2+cN5d4W2OQE5KB8d3ccxZrrjLCZnwdRitboMOj04T+Hw3sz+YVii
rUnhbj3SGEUG8uPdoqhIh34dEjulF5iW1N49ng9pO7bie7SY8WTbtMhik+EvjPq+a82dQAdropLA
8QCMyYe9uCTaSFBzI8R8w3ihS3O5FRynDdjBDDzRloytUObInKJd1Bucggwusgz9MrOP1prc2pjS
gi89gNfsc3FzEWFBiep8Pes3S9Zh13bCZ3WQk15bDEqdBoTZHUkjahk1qJix4fS0LwDXy2OY6QYs
Meh4AB7y2CYHp1RZHR2eKWvC5i1N0P3q7KvpfIGDFzpMVJsPeVvG+Wysqaf/5975cdfX2ODltvvb
MInNutPzSL4jx7fYYubZkZ7FmkOeNWqyw3L/EmdlPGXqIRDKC9vlcJyutrxKaxRGBp3mSrVifrxE
iMfq1vqFjeCN8errSuaSH0H/mHOzNIGwD48Ld60xBGj0eA8Bx8ILk/QPj4prLhAdPmMK+ttZB4Lv
/eY4L1nRyASiX6x0e+fQ7YkU9ZOy5jfvhGK5wiP8v91+Z95XI6RFAwiSRqO8hy+9HMiAjC4ov/c9
qXPDQbFuXMW5kIuSv6Xafy0TlGkz9LIbUTMFPeR20ybSWiRkb9JQGooktFgSLRSTXdgQSg/QOUr2
SMe2or9xcKKnuvk6TJ0Bv7i6yXx32yjOCBsLhqomuM5iCaZaKg8jDVthBbfHFziK/FJsMC3AdrGb
pKPzgyHWYcnB4E5voDr5nF27wPeFMSqR/MAAvDgnjHFNQgwtjWXNE7jve/hQYDVQLzipv/uoc/26
tdElnhdH+Uf/gTLUiyOlyVorCwoLH/dT2qasAr9Eq+PGaA1Rhlx+zYG8N0M31Jv8jhbgzkLbBMRZ
QdI9tNM01V2k07jMrYA3Z2wKwt4F7jUI1Pvgi1KoxiQtxmRVP5z6cKP6Apx9ZAVTzWmvKBs8ziLR
azjIQjjKtQz898H6m22EKbQDUmYUfs7RDrZsxWnlOZVaCU4ABoabzZcujq1LZp6V3+nwYaAMChKQ
uTrQLaMEAEMRsJcYXewCh3joKEN3zzGWL9K0q1ex3w4p/b23+H1nlx4ZXHpXacllBB+fpa0bzCxh
AQ/r13D0a+ndoiV4sab1HSlvML6GO0C6c5WG5lUS7cUR+usXiafZf+JUl++KU3v8kZ3cmdVyrtMC
j+0a+xzKPY+CE3tFLWS00FFy7N0w+VX17SAFrAb24DxAa7BkhQGTX/XQjG3gizKGNPhjOZClWSRA
MiKFk/m9mzKhhe9+ZIcd+wwnQKceURnkBu60vy8hBdYUoodTppDNNY0X31E1Z8ZKIteIVgy7f7YF
tXsg1YZnCeKKWsLk0cIXV1C861NfocoIXT8g35+F7WkMdsQFr08tUbv3ZwK64ydLQyOb4dKP23o2
TUrWtLP/pymL6qLvDgGoe/+I5I0nHs2wWQr6UTamEv5a9UKevCDeT8ScsFqzkZYw8HXo8//qx6hu
j30u1J9Z4kH56f8y9vsC+FRaCYO6aJLskhylzX3O4gJXRjvtdfloaZ823PjOzxVwfy3gd/VQteQS
IjGPu8EQapLE+dqyroex+54Hoxkyo6iSG7IMyAwK1iLcoagMgUKVvf1cUJr7PRUCpTB/GFoBF3Q5
GCMQHrQE/1drruAQasGZ1726SYFZIzjdG9K740gJNxfLH5vbwZI7iNsNf3E12JWJBmPH6uPGlz8I
gRHMHKyL5e8ZD2fKWUdMlWa92+SHYIIotyAfW34K7Ymoqtj5NIZH5VAV8x2SlPOnXCRPKp9lqu3I
7uG7ayPkm8g7Dqen4RbHc9ByxaYXbaUphgAM4eQeIRkuhBDaUwVjhcy0+wP9JBm493uWg4CFlSJ+
rRicKRPR8Vo8q26RVMGwbpwOYw6+T17ejiVrrrrkiqpzGoztY1sgXU3jt9P/ZtXpQhRF2vTFzA+g
gR9HVVHHC4AQHIGkPGuaqjEdXIEycmMVpflyoYpobfgYMb/hMazeqxi8ww3Fb8YNkFJrx2+tp7j0
s3r2CLxj5xai0LF1OmFyF55PgQRkygG6kYBBkUwnZbb43sxuua3Ih7GwlktZQKXeQNoe2t5LXNpX
lSGWaQxeBSDUaHyGxhCSGY5q4hKRyixY9PnaHywLrzGAK9MDn0792muTIml4VUgKJUvB+IYbIleG
CH971vmp0+1UH1ySLnRY5R0ss0lsuUxQlne0EGjtybPRPxwtYhIiGF+I3n2tKiKh1BrL0ePnXb72
9Ot4oeWwGegvRihJXcw0nShSyzaIP/BUPkCuCSjRz0UKviEx8AXgAzvnYnqq7l5DjihbdmRzlWDT
KuTS8X0XMTJ3QHNrnzHeVnvyEaTaL5UBmkNuZKrEGzBLt5V+8OPh2iOtrh1bQwcgxCpQTKOxYb1o
vrSJ+QzcT2FV/zyuoRFTR12CtxWZgDP8Wp1RhpFLP446ok+ATWXJqb/k3oPO/2CvIZE/2ugavvQv
HzeIYodGz4K9S4K3IAAkyDzXq6RJwdOxnRODjZGdOg350sRherLnj6VU3gZt3w5lnjMSu+kdd2x+
Jh3EZxvA0SDGFTOw6omKnMgJlIHcpO2xHwv6tUJTMC7VYCeHocHhEY7P5/z6ZpYvQtDrb1lPv06Z
Kblwws/UuWVL1FTMor/Xe4I/IPR8vKVq8tZJSARI2k+h1i1vU6JUHJeBvMNXltkLZWLcr/6bWlH3
rkq4mbCALs0oFZY4SRDLhWsZGfUYjq8lY/9Do/xLzWfxYFt+ZseR1+YQv34MR6PPS/BI7f3uGWoc
+T1EuYlnlNfvvnIT5C8bs8baJibkPOGXR9zs+MJWyyUjtQr/znN9McCaEvLvjxjlZso/2J7RpTUj
FEyeIj65TzPzq++pwbViOM69k/i1rdC+OIyfUwhYEzbLvsqoZOlxJkO7Z/efzX2TeyzEQ37JyFK2
6LNGWe/0PJPr8U7rvm9VbGVDeQnZbon4NU3O2/35RXm/Z6BaH5okXa4hTciFaa47NEexiuFmYbea
2KrBq0JNqCWqR6sKZIVB/CqCn2LHwyFMjyNM3hBvXvhvvuM0JFEGqFTp+ZrqWC5aOJlD02iXA8l9
aIwygidv15SeKg+DqVZm4yf7AhdQgwl2so/kh6rY1J2qrjapDHRWPa0vYhFQtKlLJPR2PPCWLYjT
FELUemvQzSpop2rb3Cb0H/pr/El4KsPhAnOEMq/InkpmPAhzTcmps7prPeJgjmGTd0u8BEoWMQkO
flJ0lsqocP/3NaAgLUuH59vZN1p4wRP0/FaJfp/Tua1BfbD1FcKQhae/1Sh/dRzHh6CdihEjbtyk
4J39GzCtZQhmlxZtRMtDe4zPkb8yMXO37R/TtEaXd4V0uAoLSRyjYqWDM55zU8sZwuGF3KXdBDAq
7K0YPpJUM9t1GzA7vRIhR2hCw3cXeVkQutx4h+y6nKL7e4E1nJfYOPoEXeaxhn9+x/CmntQA6aMu
Eh1A7/ZnWYZrp9EzskdYsMhOEK0OppgHUhf5pkRp3miulgo7LgKoDShVjuXW0HYDit2lkhw4sCQM
ahmVKuOQNkGJYslprVjrSOpMaYINbA3zmFaBI1H4jEPqx6tbpmjSmz1zltSpYHUcA7SsssS9I/C+
RJRmYPlSsCZfFkSKPyCJV0VG+Ohe5ZnXSdhSGR+XlkAzxviGl+uadVuqQyFtTzkeknfm3X1IpaSi
nQkCHalKUzMVCphlAUSb04zHe+4M4yFYg6WR9BUD4TFjLYPX7acklnOpUCb1KwluzKI9mBKaO7Fl
TUw3wTXVcUvMMY4NI7WfcGTJNJ/Lf3Azi38gORJX6y7OIDZQncQVq53/ZVPtWD0jZ7iPedSs3zIA
83c5+p7bixZ9CCE5I6+5FiHGObz5XJwp7g7eHU/3S0XvG4zrMzU2ggEPhgSvvK3O+enk1riUvRga
BHNfXlR2uLYpppERTpIjLPTFYcRugZriwnzg+2EQDRINQryux+1StDtYiInksl6VXJsK8/uRQkmW
XLv+b5ASm9b2mdW+a5QUz9HLSNt7QsWojijX/cdXTxdUOIZHlYtc0VYajtzjrf8E52pbdzg28kO4
FfNqUBumZrw6m1bY9/i3r77vh4rDF3AqOoPCknO34APTTNWJ5tNjes/ufW3Mn+mxjdbCUtUqL/Ua
13qkFckjqsuyogt4ek0ot2VhD1ink+yculsyC7FKDBVeCDAoPqTROMRA5/L4P07/B3L0CZoOwEGj
X3Hn9pOTxJtfibQw1ZvKM+IeXW2NKNhjQliagFlagBZYWyPY+QaAFAiuvLG6SdEXZ6Uk9W+tp0YT
X2nLxl7TyrdC/PCTl1Zjyxsfmhih2manVbQmS3hrqXEsvLEOkODeMbfRMsMXuZht8vu8puoDXYnK
ChwSQmS4jg7fYzJSidjLWP00nfg5UHZ+3wPNshSWSv0mqpf+sC6php1CE14T0MfiRfCeFTeqAMYl
f69Tpug4kzMPgM0R44e1kckZCcIOuxSBnz4miAq9K6VXo9Bn40sWaidLH9Xt8/yvX/k0o2HcJed8
UWqwqGolRwkTN97DaLylsYmaL0O/cyL/JW0N/DpK10y1ZwgunYuT80IydWXzUOwpDnV1UXq5QEyl
dOGW4SNdy7zhxiaZwZxMSdpAeDCa2Xv9cXpdiH8bI64RJpgghuwEZLUXcq2GQdB+j6mJH6ef2sTT
t8MVhBtT/gI9aLUViYwYB2fsIMNjgC6qN/t9HUgOxVYS4PYKWgm/RbytZ6vw/8AHVr3sWPdIPQ+D
ilEBOb2wH/qXTCE/TOWPDOj/1eMuAbtAiZnewrkJmC9y7mQF4Fn1S90kLuZ+QjcCW0qkOqys29dn
SLBaCQ4LI7qMY8UJ6flgtAWyIXzvCSO1QgZRKAs/5vC9BCdB19gAIRpp0bzTCTN1ejWU+IWQQpla
tHpxcGHjC5blhpp1N8SEoVuXC3bEOWQT9D1s6hnaSAOiW8EMWbJeOT+rxWZRrvzqe3DyyxHMiWzU
dLv18hW+sL1lcDPoHbwV0PMUv6HFUlmfYyCTR9wwJvKzzIF87fOHEJ0GKot83sEfAl2MHPbk6bIq
vUpihzeTIn0/ZAaoGuUQzVCsj+eBjKBEOCjiG1FoXxjvNWlAbsknPdLrWCfcj1kuhRflcLwbXs7a
ROaQDkVoVX3jfwvXfpFgNQbitV+18RhbfaDcORdDm0UHx6boCuezfGgwvpd1IsslBdug3jcmilNx
wRg3+o4sE5GEaTQ2uu0jhFZiR1mCvGb+jEfJMSc8Wjqtb61wxqw1tittEUpeQpWWesXaWlgUWYAO
5QNZu5re7kWTfZ53rG/ZUTmCWn4G3M9jVpFTUpU1Ok/ZYZMagjGvKl6a7qhAYZV/M9NhjQDwyo87
Q5Dg3rlxrHlSWEFJeFS8IpAB8tBgk5Qmuzym7rQqjkznoKTjrpHpO+DhPo3zDp2sQS4Hvamj/GMV
tnPWEhGiC2W3q9GIgy07OOHGkykf4yvoNojkuCyzmetShn4TpLQ4oq7wxymZrW0jX9/PLUcH4H49
bHDbJCGdaleuMK/NtxGl2h+jNW4gq9kDALXM3nV3n4OIdCKaT4O0iyxptnu3mmt0wGIeTiKS7eC6
OxQDX6EQhz4T1r3oQ3gijzz/mawfYa0qwDwI9ptZBgqR87pAKcRRXiW4M01lVhd4UOMyy5/QZflD
7K0wNG0s1WmKhxiYpG/GlCwHjo1jSYQUZZbTVdmc/JxcXReLhieW5Tf5noQahCG9DQJxRkkWBOUb
oBCkZvgiTULr48TVbxDmJVB86FUoqCYjU3QLegtdqmK2SEpwfpAvzbDaci9cxq3dXiRaXM9kA4g5
TNoBT1fuD75e/v8Epzqdbsd63rnqXjG6+Z0fsfxxlXc1OV/DfqXGjEzmzCWGTIqW4P6PmASEX+Id
RS7jTqgM9nO7TTyRVz804f28yuD7uTXsBIam5Q1xrNPrQT3JqDsvaBmrKzT/yUVLtTo9ZT/WHmoQ
D0uu303GIE7r2rD5PGf0MYrgrbswrF6einqEqE/Git7cdIKbnbTKyJNQTZMAm81wFQMtOkN8+9oH
tLV1T6y/ReJMjIFz6tkwS3Z7zYKuIaSrsFqhtaBlYuRWOOngKp4OKm4zt2gHqkbkmpNRARG4gtF9
Vd+gYt4C0uWt98Uui5oAa0Vaia8F9FVhF6w09CEMG09LgFOXBO0uTc+EgdTuUYtCF559PL7OiYmr
pdfV6l2B7W+CW8GcB394MaWy63wiSFv5GsFk52HmRhwFR8agl01sKqyDZbQYl9K7wv0Ui4JbvKl/
4d+zY0xT6Jes2NXpgBkP/ZaPMhXles2A35FDJIbGGgU3BuyRzoBRBtr7uJC6Dp8uAuhiJYuRxCR+
DWU7FzuO4zoWjL02ZREVNuWI4MewPKZjthJWbw8SJk29kHG9BN1/yKGrTTa16uvpFpn/joK0QrRq
0AwFlB0L1T1F0OIYolWxOqHmpWdJ0InsHy9AAR22Z0a8sFSCYqu05PzgFlon0HqJ8IhnNvwn1E/R
AM6k6wZT29SbuuBvs4VPSHMkMjmOvsSWlMgETut49MVjVYpvi96CG0rBQ9RmH7sJ6di48jvlN0GM
cNTqJA8g47gSYP/Qz0YKHYVh6u5g2599SSaGF5uspRF1EJML3NbiYOqxMkQwi84Pj/cOIShLVQr2
OiHtJMQkd9UrJjjHGvR7rw1ghQKNQfxuWeXKAZfQBHmLjDkras6f9KmEcLoLLotN1s34+BqxJ+ol
cUQumUMOGMmsbde1q8TrAfSlYKK3va4ggl0zd3eGHzvEwUwlQAVyJMMmjx0zraciN6S6G76WEYCA
mS165oJaQYe6SFyYq9ihMiaFjCGpc0mNlGnphYd47zviFTLzLPR5NglIvrMuI5GQcOnKpkxTVjpP
P1obxrpu3rC/pLlVME9rLB3Yh47XBIIV+z5WPrBi0CcHNGoeJuNeWzCr6hxA/c/HIux9HC3ulJhz
8IzXukOidMJIc8lrM1VRQQHrH63U8LwoolZ/vt3Z3BuIJn/f5bBnL30FD8zdakT9UAlxRaLrfQ+M
wFoiIQojkXks1mWrQgJmd1QwQsxf5qS3FcU569P53QNMuAvMy+JsCvBzNhhy85NUJLdXmbSjVase
Z/I0EOkracNvFwysJShfsmI9n0OhLk9xo4eapW/PnbMj4whtcEfZwOPh3TjFL7NjjpI3ENNY3Rfc
+RM3SGIFDP7rNav5rDl8QEgfj5gG0ByJeA1Jyr2xhs2XYDfekNd+npsEE3CS9oA90xDFRMg1+ryR
2qrvOjzipCb/9noqMNpycUqdoIXZoF1riMfPOF0RaIi1SdNnvmn19F1MylatcqeplESkrbJOP4yC
W0Jq4qoWRrCAUNJTd+i0o3miODSR2lxVklfM6VCbe5PTWMck+Z0yZfRvI3XLnKRBHcaa8FYgMPcq
mb7OGgbEEkqjkbcDH9o5gGLnHIG4I1h4qYjjgmRpl96+JRgE8TiKqRHBWKX5LT3NU0AYaJldG7cS
k1TJQH5n/Ql8MtbZwyJrP+tAo43Pd4RuZRhZNUJPSZ8XuBBMRetzR0dc5mihdu/Plli/oTXrd96V
IFljw7IsLWyQdnzuVlAW5fu9LO5kLl7Hzj9urK6AlwQQDsvbmWr2IGyVTV6qw4HxNHxps0Yjqxpg
oJvMqZFDnXpTXh27Z6HB8oAEGZPd7alQdnW5DPpUpszWTqU5/y3JXaxUvHfZ8YWXgJ4Y0H75NWXg
edN7Z+AyvlolDrddKD5nFziWonkg87v17VzpYteuc796pDqD+wnA13QdGSrdmAfja8zCDgxD2x6Q
4Xxd9AnVNrCvmJcJZeJMGi/XHwzYV1L2s0u/LDG8u4jRgcAUiDZ1H7oVszJy1yXHb9p3TQQu8C5C
cluE9dMfvIjnCAj/auA3f5+gOxPocrAGU+hwsaR8JxAHUpywY5vE+ACATaPbVij6x62FA2ND4cR6
ycRLoHlsN3pqZKvFzxR837XVJwTDHSR8oghTQmAhHqIrp6uaiAmSCV29n/EIIYvAF+H8CNn5SGiv
mM1B4gYAUxDhPFtSIyjwGkOfbD9MqQLpAD0KMdiIrVSuRgkaCxNLpnlHmCSDXdrlwcdCOdSbltP9
+KCJWnrw9xx16/T2U3Pp4ojaftp26/FA7j27ynbb652GS/6DArhRcxBi01ZjEV+N+pqWT5puFUxy
txQWzE4yjvQNoZ05t7bQ39VqZjXhMIM/gg1yfLLD6wu/AH2CwihhuViigwj9e/vYV2Gb5/hn6oTP
RSuXyxYSivR9ksI+zLA2KVP/clCTkZTOSNpvwck8xO+TP3PLeE7wLb/IrUTjDT11C2HcRteN2yAy
swcnNPAbitAo1K4LzV59yQXiaxWXIz/N4jdHt/Mftd9Lel8m9nWcVpECHs3XzJzsFiLJVF7KsPe1
HOeBnbiSIlltQ6CX7gYOXZ6U9fyLPsPh6IwbIyhmdE5Y35iFXWLYeyFuhwyjhX2yUi/Ri3MYns5R
9nt4FPN+4U/hZVdrPerZn4sEIgNB+68I1IdF/vPoIuKLOPBWO4OK9cDDszc32rNOEPFEVa1qGfib
JNvX3IScYZwiy3KyxPdix+v07iMPZ01I2qNNgG5tbGqDTPXGs5tOZ1a45O/IRCO7nFLPK1x2VyTI
82aedSaBSTjoFeY3WQSF09gX+R9xIYQx5RDyGADSq4pefffcBvyidjw29l83LMnzR9nUoMbSx5aP
tPSKU1Ogc0USJB20P1Q9gCfMzdBobj8sNxN9gidwJMeAhlanRyG4Ym1FVfrnQfUKYedduenc/G29
4tkcO4SuLlg+bjBu++2wmPL0g/tTZQl/om16XCkK+1ilvTmO3yo8+Ec7Quq9l0HS3f5Bi81hvncN
M+5qm182xYprfSj/Yn43tV86UIMN9GihdNgbjgdjkeWbpuOZcHGsmwQbmdrKZ9GZaSUr0lr1FiBJ
42BAbaMwiqhXc1p/lpRCFsy9FoqVep+B4ii9uBcjDTxD7Rp5OxUCUwtKVijNx6tXDD6Lr01UxaYu
Z7rskSDd0C72ZhlEuSY4meL26NrLDXOmYazxi119EWkFYRJSkzhZca1EE42IkaNf5hE0yAx+KNZx
OnOFRNugAlA9qVtsyc+0gM2o+Zt1YOMnWtY6gDw7akyzV5wYcpUiG4G02S04rsBVZgym/RDJnbye
EIed2phzpt0T7GsJpo4i0Q94s8Pua7xXuYVQsXDigHSafnT88J4eDGZXvfHExCHlxiQ+/1B/6ROT
K/oibbpoaazK426u+wTnM+h7O9TYnxUozTDgeRAl+PqRBAJYKTj2XjNRvf3Ha3MVU0yvn4/xXYEi
hE+Bg+74iSSOVBTVq2M3xE4DSR1MTvBZbxMfHVamn5A2RCJiE/MjT9x/+5ImTbVvLaPWb7VDDbRy
4c4yZ+O+XRgmTB3sdoP990ixfcmZyxsKwWscV619g+9duS+ueU+8ZX5dzQydudzJVZThAWxQMeWW
P51ZVcaY+GV1iIV18tz5ebTfSyS81GLUGiQHWHCXnm+vT8tB1FlcHSP2rgHuOGKg+XisM8jYTxuS
eQRsbX15pSiNJRpAC9q4XgtwWl2cnNQcoEQNwrGsi7e3JyPzY8g5KTOBxGCaORoBrjrvrcLMWcdT
SP1VYxU90NVMLSntcM4DWSsrr54IT8YFWvyUh+I8c+lgrykpdGdJr+lM90hd0UjNViSgUwjHaFQM
rAxD17Q0QkZtlxBJKOg6zvEkeF2CHr2M61xHJpeq2waXeg910PEsfNtBDt4uhoUtwJvrxfP1Arww
QLaRiB8dG72k4FP6eCyqU+xwdbj3WDxQAbSOFvNEiS0/SXpJBKMEkcaSsphVjeiaxsYGBsMNSoLl
gwZP2CUUcDADa2NriOi0/iwJBDnRZG3rtXVtcIDqGgnxl6615fSsMTRI+mIk+KIP9jqmVQHG2hK8
EVdqRkjYTsrXHS7ItWQ5yLJjvXuIwGFbrYLlzlZLrmKhdSwkGR2dIKTl/GUk+85qTV8FndIfPRCM
6IaCqOPD/4OA5cWDjZIo5oTmR+4UfvfCfE4IYTxM2y78pd/qztLsbruv4iQ9NbkF83/KoCqgKhmX
z780zCa5QVe7u6LqGbIGjFTp9aUtbavs70LFOglWJCgVzOvsXmaoLJuIQigbl1id1QxUXBFO3hNQ
0u7NQeZYqLs3dTRhr7LsLYNCLM+ulb0+P6NfPb0pyb6PGOqIq2SIJO25WuryD4aKkV2aXy29yDas
dMXToRel2PG3TCaOqQFA0f2V7KgGmgmEPJOdABMt9hBWynrXIIkwij71Whx6SfwirnXWNNwxbWf6
6/HclMSVnY5tDP6EZFOTIad7p7uBt/xyS3dyG9corU8rDa7fOCN7dxOnG3ZL6xUHraYiBwSgCWuE
eqwgz2/M+kgT+w59RG8zbrEjst8FGpZoLMyjp2M0pH6IZGQfnen6xxakWOcQYK7ns/L1xvcD7Yy4
YIFbTyuq8+72wZPEdn0qlOjkWMyqR4ooGgJ+lKOVP5pWDC+8AQ9oBZuCzHQIzlSlq5BwTYkyx/eP
J5rORFuWq6cGCCF4S0TaofqqQ/Hihhe/tA9z7ueLw3k/XPMXzgKqe4FzEa81+zAGDhZQb+M+Brzo
nCxNv9w2hZmNSGdhVXS7PP2dt1y5T5J3jax/d5SvFEE8/tX6MxW2D3ODDlNJXedroBJi3Hl9mAcH
KBVCdj0tRRng9j6ocmkU+8hHlSpnz8C8ZfxtAwl3hnfbJNI208z/CRnL+yqb0Y3dhkfSEuSv/5fF
nrdswrlC0Pew7JyMRdUVPbhUvhF2Ofq+9cHLOxWo4AqvT1vmJ9Hi7uwZggJAf2wkZnJ0m3diAWlJ
nGeCpzcj7g1Wpf9xtfvJye8WyQfdo2ZFqJ2WziUABUFKpri8EIT6EY8t9jpyaj4fCNXKsPrLjJDU
524fi7/Ilw0YSdM66cZAyVb7GbhdZdlkbKuS/DhE07Mc+WoUlK6uRxjXk8t5ealoiS8zpa0XXixi
s/SM0f+Oq9VSksdBdEzzU80XVhJzQ+xbd/vLfRExpOeoFnisRKXXIMAaJWnAJt341Rd4yduC+9xR
xKZfmjY50S0/00BXjJkX2GImzD2mZBAiTRpgBlVscx/CmEsxs66maWEksyWL1OAW4yddWnky3vb6
/Apa24Zp2zlLWm799R2t4ub0WPha5y2M+jqorA8WL1cIbCJQqKkY/HtxQX7AF0CtsKTdWoo2n2Nb
zCfSJv3Q72Wz2HacsDhe2neADQyRV7vgBDtU7HqMG2HeYyVR1vAl86i1lgXH3feFHQZhkQ4AkhWf
sG6Fet1GiUpdyfmf1CmosZYgdEQ2KkE5dHMQ+/9ovBS9EblXCBDVPbOEHxJDyfISNpoJevErv7tj
dqY8EZxRS033tiZq9SVyiDgtlB9W8o/XCSV5WkeHVMw7lw8wCjUgDaF/f6vu4F1dBNe22wWnFMrS
X+WDTsMqGZVknR82pb2BgM4aGSIfHtayDXGi96ovgyRFLDw71QFFH1ZY1BsZlWcqA7X5q0ZmwBFO
WftLykZfQRUyJ71lL0ZfplEeIhQQ4RQtbjswAe8eX3ntpg31QkYsv7bhC9LP8qoI8k5V4gBN3KDz
m7R4o1A5jKh5bS3CW09AK5idFWTMK5tFFOzV8jphVHsd5fg1WU8DHBtnXTuiwN+q47eMvJabuyqi
syTDEK/eWad9Dj8vih+qbrgYAH1T4cmgSSBnvzqDolMSh8b12remE5qpo6RlR7jKOz2D4sr5JMcB
mx/l0YqGH5ycXKpGobA3YTnhQHbFYsUu8JelrS6df7QnKqpf0IzfqbIIoGsihXzVU3ytKUh03A5N
6xkQ8sRt+thamnj/vLNgN2j6def/37KyByPzTCacjGjR+IzcDvGp2UX3qwgMDhU7Aeiyf5+Bhm0L
fty85TksEl2zVVEz4dTeYGv0Ru+3IuaEdDC0U4FK/SYmJZIwXAi9BIOSlNuyX9C9JYXduaODVM18
XMsjFrHjMdGkITJjLeWyDgsiq+vGaUc2rNxQbf3efoBaddMSkw8hHOkAGc98VM5LTROnks4PHs2Y
Eo35OeZa7Sx/NM/06Q5+LZH+Nfs68MykhP5fJ/gBvvRotzw0e9DqZ91LvfvhMNjLcJvjHRxBMPVv
t4z7eeBgF4w8eO0EcLRaTcyce0vzlbJuXBw2YH++IdetEDG0ltqOxBkNPEe1M0515hWu5ykUIDUp
ZamzzCXhbKBTS+q5GBlQhUPa4yr5fixeVBfs47L1L6jNQfcoEICsnTBA2N7fM9RGBa0PvbczpkYI
da5JG6+tW4eiW1bKxrS3+N0DcRgN1XBTedH0Ghb81lIBhjtzRPJ4bQ7/hYZ/UfB2kkMsIiZpo2WZ
L1WAdUOEco4Z3L1vjEZPbIbF0e0Ne7CV9Mmk6FrJCCsJTWw9yvtP81kT0wBGcWgp+8ZSuFAUeKSq
d5aIaOCNBJXZgO9mVfS3V7v0m/GoWnP4KobxBsa1TM0kbjkX8CoC1PvI4sChGFH4Er4rTwAXukdh
SQ3upDXkmWEnEF+BIT8A7v7hks9CdgdORmHSYOrC6lz+1XRmBoHVmQTWZfChEIELk8k+dgZH+4lq
uFX7sAz99beEEQNnn3gK2C8UydUrNBYBIybqs6jD722oiViKyAnVFBB1iMYM0zS4oT+G9ic3eEYH
Ls1mSHaw7G5V1cGIrI5ctI+Yxm5YkFSL9PlqdJyluuuWUuFBxUM+ea+CdDTozw2vR0tvIADQGdTa
U9K2zjHTEyIS+TmsnIK2htmH0Al+pg+bV0qtuYt08sdZBkHW8pgXRVTKsSsQkNnKpVf2hbo0Inia
jXbUWcpUs/WQnx7iwQ2/rIeJsm/iGjK9GKgXdWT3LpcevyHLtrcOayzh7LDl/npYjy/jjb2zlCsP
3i+zqDwmjqkLWi/3gv9cDZEodEpxXa2bAL7ELJWqF25iUnrtWqf8K4ali0XpCavhRhJDVUqhcS9Y
dtLGQUCWs+GdGT6F7H1zn3DNPtZkx6ntoCX2MlKAou47nSoIG2/3qvZsnUK6pfE7IEptwLmoKLzj
ZPqwDH1tdr1tUNoG/dWk8wqmkJd2TznKsh+zpfRtIuSlRyD2oksTTDvZ7i8y58IP5T1jOwbYaMo8
y3EbjoZarjJEpnSQg1KtvFE69C6xy5fSDGmyKhxFJT8z/WKcOFLrLmLryeZ/ZL6zJvwo4PU9wdsG
i59sTnXwqAYzLHWgmKl1ye/nIUJg6284/vxSxwliCqQvyGDfkcTy425rWIs3Q4nexCYb3N/oYDlX
F3c2Ny4VzTqaVrTBPQNqcFYz1Xdm9Onsvmlp9oIh0YSFjDhGHfHq8NM83HSGnhCSXX6ZTy3uqg/b
+rbn+JI9r4QTtd/R2awx59Din2cmtlOEgHBvfZqgxuIFsQscO40nLhtI60kibwt+hXkDC6iz1ZTq
7mo79p1DZ+gp1jrXfSIz6733JLPYJeTiaXJyRj89cKnt0pyQyf5tNVS/WFN2gPK4FsZk/0E6PUmD
lZXcFdjj4dRJO1ixbBwFOqx8ON5tm8veJ3SFJKrrI6RlzRGe2d59HEF8Yz8XjVUuYONrOV7R1gCb
hiR3nIScv4s6ZwL0zA4DoZSAo5ZRY4t5MOkhdBqqwyk8RGXyx6In4LiYjFmilARa64VRw4pWmc8O
hEfGmK63QLFB3OHIba51VN40SjlPARbZRcn4XYMN9lQniG04+14kqF0YHW/+QbQyyzj1M9SUaUH/
BRZxOmTvJ3QHZlKqGth/F01XOdWXUfHDdLs3IQc4zIce/r21kDEt22lKATUDjFgYYqNQqejhKJgv
Tq9k5OcjMLvgcApNojavRVAJqaXW60v4kHaWaKJG6bZ9Qvd4wsNkmYdo1mXMMbROMQqMJkR2xLw6
8rcJVf3ClKs+xuqvp8czfpEpHKB1OPzPaGm131QN4zSTY1chEzAmuaeelKOtMgQ5hgL5uzEWNFjJ
kvNsLnXCQ6qUHA+qtPk9cGJfQRG8TU9cvoLrZkyIaXRQSIWHwxWq2ajVGT+GeYvxJx/HUOrDAX1g
lb+CLS2wtcmc2Bzli3Hsq6/GDYKc/JZbFvyOx9235BxKHaTZEZbzsqF93qHIB85a4R79qryV5KN5
cawWv3qTt4CBXJe2KV8r32K6BJ/djd/vXK4OTAOPCPh6i/6R5sm3ptL+3XN2P7kPU+pGQ96QtKPC
2ARPEin90P4Twyl50+g+ofyXYC+1eAwoXiSOnCfCjPQvQaSoae4cfuzwRZnojk/Ksuu/2Upxsrdn
hLqPu0aJaNzZ/9wuY3qJ6Niyy3l6z/xWjeJXZG2Vo2YpLLTNlqdvJTrj8MMQkANKbiw/j4sDxkJz
V0SAmJIjhCBGh353fMAjvnofVjSPSAwf7alIq4vkX91AQE8g6cGG7PpEOnXnf/QfOCnrGttRgrlA
DgWbTDD8GEw8rvVjMNfj9olxmVSNNdHOUC7XWD5DeDAr5kTwIk6lNcaUq80JacfiHYM3RBmvlo09
KpqWEuvm8aLNHtHixdOTsO9y8HZsZoS8wiCMJ+V81QD8uVS7MtV+LqIRNvbtmz8kWYPq86lf0yin
Di4Abf0XMksdy/geHxFKvuM8sUzFg81WLBJ3HCTl2DIfuNGNZ/WoEDSG8nQTVxu4+xtgNTiq0D86
SgSV/ESdKdlrBV0d0jaTnhMZHI+/p2jcnGZZO3Jwmh+pmH6wsmnFo3i7H0HFBoQ0SInBvKzI+5nn
IR2K5IjHQIWVWbtudsVEYd+9um432DBegKkrrspVfJLd2V/AXc+6FYEgjmkXgEyhRjLufOpdQYpt
XYqt4MmVDj/nr72Yht23xwJo7AJge0EIpkUUZSgwSn5uZoU1LiH8sSEaL2Y74LyvUlntIgulTwNv
V1G0+J8QXIpRe37TlHqLMD5jGpqlD4n/Abw4TmSSyxoQQpYZwHP4pJi8UIhIAUsvJX4jwEAxBN5K
/ab73ieZ81bsAfe8iiAvjRd3oqqpN+GIwSYTNsiaTUH1v4DfMzIGXBFhRTVJW/fWTxulNM1U2RPM
2DnSrCGN1Ebv6+aQA69/AU2ypxxHXx9mXbhJcHKdX5KDmAnYehn7iDuAm7672NIIRHEa1SmGQoQA
8zZNfnWX795v2AyaTPjdgvSCpN1WCw5mASaUetS/WG/A/Zue+86fNQV7UayT9+VXQs7lt0oGlaJA
Bm+M1dOr3Ty3QAtrKZHbOvRCuRLBLuchWxkr9qayyPke4SWCeSbIJmZnm1qFyb/IJt5K5Ne3GQCz
lkLRBSvn3aIWP3cKAM34N9kp46LjUrxY4hJg4Pmzaze9X8W3K1jpRW/0GCDqFtnwIjtnJ9Fwuvmz
PoHK7bGBIW3xVI/pMolOATCKZ7Kw1+dYZKdLTNAAy9486D6/6nN/xOpXFKbszKl48U4GZCijYdqh
ecpdt/ef9nJQGQKh+dSNnzINfDxLG3nsbN4IAIeLgzj6/eV4H29HJocQwx5iEqeFsL/fX2avw8mu
DFppKkB9+JMdsl/7+qJ0/0fIzCAHGfS1DRqFjL8f7vUOF8bXRxmWVRVYbnMD7q9BN0aqr/gwpdIV
+LfRbHNxwGky3Rd9ctWQSmoSWNDFHWJ0g3WMLJI9710yUSbceQYB2XSKehOfvVuD8JDUM8XRUi39
i1WYLdeyHkCiFVlYmi0IzlBYZk6HemsZb/VhAS7wMON+EkhKF4XvHBk8I6805nBkVA+yJC/QxSHT
z3bV/bbjMutnjtOKYzM3nMmyqWL5ZXbh+ylKGKCC0j7nlzfrUteLYOjEl2gH3hV9P7VCocgJGTmA
VWVlsD3saoQDz8Xp0ETdhlGcDpb9P1DJCOJgYV0PKj4/foZ0CzTEI5zmsy9FZITOr3qUlzgMPA49
lFc5R4QPEpOfryuR61uKyN/gTbegOUKAzv5sP63JpAsfkQ4BuOGJLIGXlc/VTL6TUE0K7oLr9RVN
9PwbG61kd7FMMPYgGaUMJIDOGN5dg5EC4UNuFlt/ahWGtvSP+8MTBQkDZ8FZzdHysvUhTIxjfmVq
tLggQhuYi5xGJVmicddI+3Z8Nj3KgIEVB0I2jr/BZrkdK33yjA405bRHYsMXwSQQte81KtOK7+w3
pxW/2Xu33SXKp17dmrE6FaNL/rU5vkso79z5c14XfKZL0TDhLKvWnFeIGHV54n3SQj4feiDaFzpV
vTUYbx/A6ihMXI0MGVLtdYIRYVnw8FaBloYRa9FLUxxIW4F9/FNy4X2ucQR88FM9zcUCTRn/rbmk
aDbsTzwNtjE9vZwAcuSyQog9e+h6NFR3eS4EL34/i9atDshuJ+mNPz8pfOpUAJx+PjxrcQG9/k9F
YSMZZU1D2CO637mITYZg8Usd/ZRUNSGMeghdWIuHs1CdmQY9HhgBXe3BQbqDwCWBqDyGSScc3hWK
8ifcuRlG55vfYK3EiQzMpzyBHFmV9TYNWNIuXVEPEjDEK5cyixpfNkIFpZoB7eSTKJ/c+nN8SdB1
H1ZGkkFqZbeO+g3FpGpEIbrW9MzGEj2ltucIzUm8cMYEJd+WeRZkb2aPTT6I8amPm3aNyolsKOWM
xddlf2gP4PYIu2DA7igg1YlxXRQPxQQ/kr/biwMcI5oCM52zCKLSBi+acE5t1caird6a0rvmpM+P
SNhr/59gTG09kT7+mMnKNcfwS4HnKxi++tue66thXZOlirV86voT68B3EGJfKSj/F3zSYWbChkQy
gm/N8DhwPOWcL84KIzolSYqA8ng+7es+fjcjvUja1cIBb5DAV923JJpgF1cqYBuewdamArgb1RZu
1FZmyYTHzraFeNGAiwpHDmPupFgVnJ6+RO+0YxIFwS+8g7H0yflG8msN6FcK48S+yNtkvqxSqpVi
3BQFsJQp/5jzTEfZicXuVXuxunpXOjTuTLY0OQSutET2QbKaNpnmASxMBmgj6B4AtrTKfjugHTgG
8NUDbQoLukq61MgyaBbGaBy0omWCtDmlz52srDX0djsedr5MMopkiK5Zky6JgJnDCd/3omt1iTNE
w5Yh0TyDSMwImO8o63N+SYWv5/qXKE7UBR0EklTnTGKTKj7B4zIgeQF1rcyZZ9Jte8IZhAXqjqCz
0ODR/+cEhpb5BskD4CeaFtblJldVAu+JVhoRWkyV4tirF+9au0Y2kT0EStMKYJGcOfV04acS26jo
xG87RIGAQG0o+SlFGz00gnKCdsA2gZ0GtXSA3AeB+wy4vG9pkLXcWq9JbcKC4o1sM7ud5pL13Sj1
daT4E7OYRIYvxgtK73l0lp/VoxpLLFoSBiVY1w8RhDec0URYhTRDRBGR9DOvmqQftcBsREce5lJ4
R2/zqQe3t7Ytj6dHS91JZKZzvILpL2IGv/iH9LNPSerHYb6PEIpi9LGhKqEaL/tFSIkdRiWkZ1QV
NFezR5Mw/1d/k4IkU5AezB4CMwq7TIcJOsbaAGzQregZMkPpnStBZ5SLKgHDzQ5pQe83ncA8sAWG
i3uQhs+6fKV4SjFrS2e3OoHkmhfNfbiqGXZfhfOUZs2c4Coq9Ug0mNysBOviee6APfms3W3dtCzG
YXe0/l3s4llIm+w1SFQoBlmTNGUUlvbl1ht93b4zUB34uDmy5xMO+0omvKheLkBz9OS84KJUtWh8
8BtVabYVfyPT0FMtmUwVDuOGdTUvVBjcS0vpBNDtQvLQsFqB7SMRgqJMwcVK8Bv9q0KD00lwS4g9
GsN0cpvi7ZAKxNcAQadErOJ/w/IALGLFmL2buErXhbpBSfbhSWVqOKtAUasADXOrEn9VLfIk1x4d
iF50LuoubO071RB9vReoABwKV1xBPcEaNCCS04tOkxW4rKJJHK/L3oTVFFlDGxULndkwAAjg+VRi
lLgEoxqZY/lzcq7uOM4vcQuNbmpULzEeoXzaKZLeYP1o9sCcxQDreo3rlIP7ANWzXxtK4rEty1Nh
nd/iBONM1O1dZd9cBHYbGjY7sM8pygGzNGs6L8Z9SF8oW6frDfutE+BoSIYrzpHieqEO/COmaNvT
jAtU9GCsBy6KlSEG56favjJh4FZm23IjwRHVh+j/K0a4NHBCAtTV5G5w96rYTC26aFLet+w/E6nL
fj1eyPOmdXMTp/i1uJg21TOlvG+GneE7XaAU3UU0ZelZ/k2AAKJq+iyEgTPFxVVYDJTP1zUFnYQo
TIseUHm6I/dMqqlq4mI+fIhvHrspApRdCHdrz/4YXU1woeuTqPVeoGoBZ7EzaWWHC9PekrxR1zRg
ex2fXO7+kTecrdXsRx4XyfxUWNSw0f0TBMCUs69nH2YlI66F5vZksKruJYQSjJJIurEcCvlmqgmm
FEuIpeQYpEba120cWh78982ZmHFyjJILCB+W/5SAgROS/xCcTYd2r08NbimsbI4dmZOuaodbym+t
CiIPht75CP8vWj5FpAC5+yhuQqF5mk0esLh2Obd33CjXkyECOiygsPQ8LGw09Jx9xNB4NpmrykyN
JgOcd8nAe9hMi+SG5T2qiu04QjQEK54SAj6uMpNBq3jtZt69BXrlAi1jlfoZA8utPBcHphbho3SP
YQpyq6/eZ+JCKEMAW48pPjwj8H57WCqRSPU4MJK7AF3wCinaXSyMnRL3M1++37X2MPQzR/53qYw/
RXKzHVIgFIqdq7eIaUIH5HrkwB4frf3vtJBN8QqnnKr+2PIuUnrL2nv40Uswo62IHQW8AW1g0qoV
Xzos+p/+sIVicn1cxXvdPLfFocqwq/rZSovB4ZwUUpAULFQVy/DxL+c8/xYIMbRGdOy7ughc48wv
ULigkD7Ru3QCFm7ZHqh5feVC7Odk9WJDhrwWnymIR/b8LLYPtHYgZRvwRZWWosB+4o5/cAHWxlQs
ytXXPTWq8fkiuddctk03dXRg5u7Ar8O2/kVgi5SuggIobOgBf94vloVkOoCTh9AmlJygYNt26Kfs
jSlTRkyjBmWj5hj0OSYSE+f8TRjtu2k1UANFwodxsUnZJLyYmOGvaLwGRDnuG6cutZFie8L/6bCF
Rviw4YdtsxL1cSH939Hl7IifE4sY6h7H/4DMfBDST1PeHot8mGTChtycHg70Bhw2CSboy3IvDIBF
DNKYRvGGxzMVy5bjY33ttjCdn/JkAz9hCVJsg+ZEEZcru5O41kncE2P+S22I0upf60Q16ytLSYC/
QvQyqqAdS1QBVMOmp/Z5S+poOKSRyJi6enGbdwJuLGkcB0nH2uaFdfFH38boXAA6bfkWkl0Tk+yJ
U0S5IL6H4IRrf+UYNcOW81rln8HhduX0x1PuYKA95eLFSlBnX4yxvTFisFjHE3INjxhzTKVeWEzw
2/QEy8MLrk3RfIe2Hj/vW9UC7z4NXzm3yfqQUx5iGvLVmDFsq14q3/ynoz3PAYrRQ+VN8C546RmL
LzkSf+pNF5t+GKBKSeuKArJQPcxstuQfnRJ9Nh7mQ4muCjbwfxLlX5ySpZ90+EIQykmN1WeXaPg+
kAveJt2Q5YHTcgVzXtXsDBy8r//Kv2jpYGhMJGBbAlVYD1ypWiyYufjwjvl6sIdTKFNLs2c32hXc
emoGSS344azM67KU+QGW8hgbJJAHZMQKQLeHRjhbz+kDk5lCVeEw2BXptRIyw2GHZ58o7WOrAlyL
r1adKSa86Cbco7FBfCt9YmOPq+xRxs4Yilzj13KJuc472O5z1uzrVXQV5qo/0lPvFEWxCBOsOQvi
xV8qW5dV58ELl5XHc4xuv/2/JL9ELMIsZjPjlSmvv+XQ000e2VhWHLZydKqHlJO67/DBjiS/t1je
JwSzcBhosk5BajfddLyg6IfTwqZn4AdQz0i8r3kEFQIfL5cP+eq4UChz24XT5Ym1qE1HEA5SmZ+g
u52/bxaxuyDnZrHfJXYAnvI7dfAv+VdU4Ym4Gcf4eKo0gmIyZlvh5mfxuHHiBUKf9eDPh0EnKVG6
EntIk4ihbslCihypDVqRMSxb4GigQXX6XxOUnWQ4hSrYD0tj9Rq0qq5259MFuAXkF5fn1Ggft6un
pXO2fBGv9lbw3YcwpSsg7XfBBICOY/h9bYZ1uAAfS1KtiqBt7FYRfwR31WXysIXc4RDcx2LWqN5e
uOg6xGb4544rmE+rfB/sUggKlffuF8I6clR5rT5Mvokz/kJXGqEgWbieiBDh7VZQdOSy/6ZvVx08
e1N2ySPnFkJZHQz2ZbGOcx8PkSLcAIIz3D2ulWOz/QixwGPpVAmtN3/U49As4CoNZlCl/x3l8UTT
ZqzVei9jam9w7GUGCFVVrRhL3aEQ+baUkJCY/V3GmIilqWJv2JbPRZigyMqIIq4RHJBx+HJsd2yP
bnIFJzHKtGQXQq33wxDsHIlEPbB3u+B2Lh4A0Swun0Ed50u5EVmCjvvXYvRmn/m1Ws3CSFZPiHMR
qjF6LbI73RjD3vEgC1Hx2i6h45+khtaQgu+ASWgYWe3THd2/uZx/vUdXCYc2PzkfdHveZMg8geva
K6WGeKsmI6oLeAOhTTqjaIkuT1uPvqf9AM10mpU1t+DSRCY/LkYbqr+VZXJXtA7pXVJELEK3JuId
9AU++rHodQCaGCBuQrSvauuGUGMLpQ+n+cd3THAVOnRVOO1TDv2GZFxOScFPezxaNvXtJDecmv93
HgOuizoJ3a12wBLfGhq2iHjyS6nAflb9P/nhFmZ0b0RnsipNuvBNqcedELSZVxHI2fMXPDGjUYyv
GGqH4Hk+fU6X+Wua4mlo/DfvWqIQvpOqH2E7CnhP88QmyndwZCzaZdtlgBcoi7woPvjp1XD4baUy
09SvHbP+l6cIW7aggZev1SsxX9mUJL4V0I/ynX2Uu1/HA+yuPH8Ql1dpu327bDd8JfVrrQ/3W6e1
rqt9gf4q1CrsX37NlmV5FyskotYvGfghQS+zrdRU8VqRoi981wv2MXYpa/R/7qm+ZjugW97qwQk3
43+VfDAXSEDO9p6ARUA2ij2OFBg+1vHUgTAGDCuMW/c6+fm6LfUqJ0znL/JGLWVf01pOk+C/l1R8
sKC5gyunWzl4h45ngXJmNyjYWuDu5BZC1wdvKy+kHW6L80ntHULpZXGYPemAq09PF2a3igwyPrak
oySqq0Nxni+ZeSoRm8y65BB2N1xnWBL2CfQSuzYhv2Td5A/KTB2JonPDc94cjqtBSRXCGhX1HITW
//5kjlfwMQHir6/qd9WguAbB/5ES+x81La5o+EJ0EUGdg+J0vb7Fqo87CCUzcCIL5NQ7ueXFn6+e
SXSKpwv4oFalC8KnRmX0lhT+G8Vk+ONdxf6YdMawuUDj5ycjZakjdrrx/nl61AqmiBQYShIwEdTJ
smThdV5Wnnw++hXnHt/vFIQh+wQiDN94LPkEq1K+A0qD9FyJWe7wX910FA5u6iiHa1D3Z6Ubc5NQ
2uKePWbwpUAlampirSrUwodpfZQOFh5GV1xXNgknDVNH/1LQ+TGRvmb8vT/Hx9zgZHeWFA6NJtae
VaoRKckQhLDrQA7Xeuwc24+ioCfLfVExwNjaMF8y6O/y4t8udY0Qsk64jW6JhbwXbSM8gz1GDy6b
cVyK8k/ldjjeV3dpvrfTOL6OUC2p1EjApQBnnyFm+c/XuGlyX7eRvercC/Q6NtinLdqvR6sa5wOR
LkAPHXH2MaSA1ogMCRZ1JkpcaFLnwn8/48+kk/0aFfHsaF484hef4vEuwcRAjXLAXeV1y87A099v
FzL1jhoLkk3Fc2ltBKp6M+VRbj7FGuuaQkf842kX7lO+TxVmkE5NvKS30oPangfH4Tekg6bufry6
q1WssTTA9eq6bib0ZG1GtN5+pB7+/d7dmTln5daDbPUCV6eXyoCbbFYZCsy1JlXBbUIeYtkVqnwc
2SxhBWsa8uwmMVt9jpPm6g2d5+XX18n5NnKKQdEQ5at3/kBz+EZl2URWGmK2EH3uGe2dRVeUSVqr
knIjrXDybAMVqLd7rOG2rZUlZhua4GgLWBJSYt6Aodp63fky9Bl7h3yN8mcg5CKOXyegquusvZnH
/El/Nn2JX0pLkMQscBzqz+TF5QhYaNWr++p1V2/bNrdPP1atPJ4ZVOGMcoMWC8ipfR6YwntJZaTx
OT0Hxb1M7sgfiUHjCy3yxgJ40OL/R2fYDwb+Q0xxWBbNYh+YgWOpQzTdcVlfSEmaIJ6/Q/nMrZp2
Xggj31B07F7+rJf2jMO0j//YBaiNxTTs8VNqoR+0c751kItcZ+rgL7kxraMLJnyLDtPdr5jO9IH/
O2KDniqdfvgj08+kSfPq12TZltHVlA8hH77cPRaXHyLEAddGWy9xsjeBz018HcOte2ZwgIVXnfth
9snAZCaZ3RXy5LW3GHXPgn/VtmdYQR4AzOKHGh88ewPLruIIo6AE8UdiTqWfAIzwnEMAKhQzDuPv
PBKzsdkxqhZjB6KczrI+FivZ3wtGCJY1RLMAEwjxHSJB0ZGoB1pa4EFG9KPyVqqwSj71+/XwNjNj
qs5RSSpjToP7TIR0VcPtMrcgAe2I5/4deBmr3D5xzSRuNABSg3BkGJQb3U5yM9YEDNR2ymVKLzkb
Kk5PjMYe11Wzkco+YeFFlYIj8jBOaFNK8RwtyTV0tGx6r8YMtw4IO8g//8Gr+KBf4cF41VkZnf2F
z1a0l+gRgOS7zwiYWEUdfRtR6VCiUcEEVjPucaLbIZOwHVp93yVUpzOCB3cBzSFhNlm4iQ6IsGnA
WGgXRNvkh8KaC5JhOyTK13cU5IOVGkyJoXeTku2amlvyAb0SPo60J1YjaYzEBrqO6sGT4dEjk2G6
d84rD5ogqQdsiGfQ1INww1T6lVYjDJhRhHEOwc1qhQYoI+KJ3S3vabLTRR+2FDuhncDYFWydGbxU
DahrJ3kPQs98HORnhvakTQKdmEByh00Tg8bTgKCUKzXJYuD4WO41w1eKu16r4X+dlx6d/P4dB9TP
AEqtiT3iTwbakQnCArKWIdJNloy6d8sSv1/9Xd1DSgSITj2G43vFoaBmAsSLqkNnzAQGMKqxCmAY
TBPO9AGUvGZos/JRGs8ENyuNViqWdUEbCjlVyhcO4mXDkM+ZcbmpJ/N+GZuaVU2Yjlxv4kcq4kkZ
/zh5dVM8g3b1Cr0mJDBsx63Lhym9uBP+8eR+fR8+lWxu+RuvZyl1b4wIgnKumMZUC36ypf3jNYdL
zvF6T/k+DjrzBgVs3zAABZLTZ0hx9hw/q1Ot+r36kIzAHteJUiJg/ElfxH0L4yDwt6KTkxK4fvF+
7jx+NiQGCkdKeUTv1yB+S60Xh17LfBjqXiF0Z4okhqto0oHq7vG0yhfb3xwBaVMCnOPT2sqKu1Wv
ztikwy4q+5fEcm+NKFQ1ttJwRss9UyLV5w/KpBR0Go0m4rXX1qZweav08H/zKzhWcj7rM7UNCPxH
AQOiV91mqqbwOUJJbWYP++fsyhyMVmFTUvCZs8AGyCj6+V1WdmrqZNbtPSdA6W9bNocFJ4ayRFWY
MvnqPHSKFu1A2eWT7zU7SYOIx1d2bojivwpvb01BFGcFHj1inikK5fnGkSWea+aF8AWfFS+YKC+1
XTeDCfJhUha3WGatAntQhSlQRQTwzA5mAXj9lc7VDzC14gqlIdZo1xiT5B0pxSe4LufD9disiu01
t/5nnWAcsg71vRDnSkfLJmZSKj2+OBjI11C/Zelpj32dSn90zku9gU0dA8ZlUmgxKP8GSuDCpL94
4ReZ26rB4Z6S7fahp5Iud1vS75g8R39r4rLLnHg99mc+NdNXCHqgq5FhOdGIQmKS/tLJTp+zEmg6
fZvFNs0rXJVKShmmxkpORRLQH16eMEZkdadLJrtGJOH6FxBt1Ya8WRyR9ZStqJB60Snp7kEdA2QG
1W2yIeQA+/jkcHSD9FT5PLGPZ8FU32QiC/fXE3v1CYXWfjXX6RQk09IDaXPp2txP/ISwYBviR6Kd
exdcbgxkwYocA/53d8utiNenl8r7bz1ZG4x7FMPi3zQcf/Drjj7Ja6OKBCCad+O/rssSHI0Md14J
8nll+WOC2lHqd3656Nh8+v9uls/SwUFk1RmHyJLZ4lkktSNuFt8oozmgQvctQOl9ETSn6s7APQfW
bC2n4qEZoyry7tv+zS4/u1sdNU0EAP5ewDf6Ocpe8LfMwjiWiJ13VTo+bWNfLuODwGdkVPXACBKJ
zEweyJzcOzqpld5ROXXqIGGuOk0IaN0EkCJniLV0ByKlWSs4kDxm8haoplMpT8IKM7a50QDFhjPc
0TDEKAVUcCXqjd1INQALj4mw97v2Z7jqMNtt58OK3hkcLLvNlLGOXj6uTuX1y/WAOkO46OLK8CQs
CYCGP2LBiByP+GZ6jtefrJbaxIr8EMuNJtNKhJHVaRUhgyUuxkf6pRDv4QBlkMGxS631GEB8bcWe
afG+pd+d1trLV5uNjsba7CuhFNwGFzKZgc/OcXUOJ+XTATG5+h2dw6GBMpEcqfJAEs5xQv7w9qCl
a5sjujLINzDku/eWX3Y6E/ay/oDhaPw5VGZ3tui4jh7S2Z8wMFa2vFYYmIO8Ex6w2ABIfFd9dzeR
4M4+upkoqFC3NnUbBAfyigGwK+NDyMPeB3QFnPgcwpGRg9FuncGEqcWHN4aWeXwgtJKTsVw7cjwD
eD0B8IEcyXpcfWJG9ZemF43Y3NRLOIywi/9g+Po838v+FolWL6T0TdPVCQ62gL7d0XpxBh8hzofd
6uGh15iZWY3Mc2hUvhaLnVuhf9Df/DG/yrhRCGpfAerPZPGD8wfIfJNBcupuSv/MTByYjZAD9+Ze
Do7V1Qfvlq7rIK92smSwPlgEdsgVL2uhpEcifQ3U+VWd8H8le9T52CQiox5Ck9D98Hb/Fd3GOuuu
aXdMacbvgtojM0Uj9/ax1PnfCPo8HZszfbbPiOia8BT01G1wVB33blMN4Zxdvjj5pMbBVFdvWOKB
w2Pa9Mm+a5DbeM36tEkh+Ru2sNOuVB5Zgajsy4lwEfCSSAVOqZYsoLgkIaVRw2UlRIQa0KqnYZjw
UuMeQDJ4IIj1aBMSHlcEQNUEqz4vmrHrG010Wmn42FzbGp3lMVsEqCTWBhGiSHkVCTRwEwPOt569
WeBRSyujpWkDZpcaM2L0102VgbLgBt6fSOeP3+Z65SUiJ4OqP8WJRmQEblHzYv+iA7kPu6An2++I
fvoB2PrgtV5mla3z+cUI4NPWruCSS5a1USw0e1EsIjeLCHp8moQ1lJph749P652twY5XTSVPe5Jo
a4LX4Mz9MHAVKGnxA/owAzAsw3gt83O+Qn3nckecDUx4YvaSSVWuoNbNOl8l/VuaVBZD6a3Ps3rl
WXS4yjgF2NAXJzX9v9lBkAtKCnaOoiiZrBRQhzvCXKNCCVE5s5Nf0fJ7zB55hrtlTMaFxqbc88ET
G7V8+wTRSyMdInh2bQCUhZQUdo+J2HmyqAoNccljvNhXYazJzLFiQ+Mb9tIkxqzB1JM0sPpAMUdf
emH+quXdVVEL5trZWvQhNgrQMqVNMPQSpozTTQfZ7MvhTBQ2Y9jvsnlfFy5AGPvvKFN+LfGBYe0F
Wvk/wv3NP7FRXBUnTYYiWV0fgH0WFMBEObhB/vsoiR2e4W3N4QdpoyImTF0vWvyuDuuB5esYlzJ4
/egh4lPEIml2fh5K3PAs9SzRQtrCMlz+s2wSV/cGuO67OHtg/XPH9XDrsjTmbj6Ttco4O9iKhiP9
k+G7lq44IMAxpOezFU5GurSgJXixHKmP/jWTsMxKGrHoMzwSJaJfrzFueg7illrhwDqAE7m47tob
x002TxrzZgA2NbFmTk7pwByvvuwjRDlCTJl1pBMWTqqcPYVDvrcz2GFJ4oyDVN+0tmZDgWaLCZwy
UOR+K99NGNitUpBP7QkXQe43tFZFFTPbxjMp4sluncayUDYwV8qC7I3+cKcjFXtG830+d4sj0SVc
zbpHRTDCPIpRLyNjQh6D/xm47ibTOBbmQcUqz9Wry3oCfg6g5r+5a3L/LDB5rkh9QI10UX6HNsoD
o5K61UH5wrc8X5zOCOsHc1BsuOOBksocshDKhbmIlyTHNgImuhXYMCfB7IgxnmOHhpi8PSq/w49s
RnugG5MsCATtX4SLr6ZAKtFS7TH5uOEc/WtBOTsTCKL5aU9nTeEQcLpD2C/wGurOQdamlPBFRL/7
vJdB7SqH2PMjwvCkqbdnM24x7fqhOYJeIqjbmOWRn6027ZI714XWRl/zYh6PItRXFYzoDPk43aEk
vlWsnuINMazvUQmop/OtvJZbfKbHtfKbN2jT6O9HVta9NqkqNXRvGdUPiisHvM4stSUzlU2t5wri
87Nkc3iAql4x65yFsTFWsMVqzy68kQAPq4EtyxE4RmJbpRYSbmcMuw9qRdag2B1HR/FPmwMJmBhC
gwx2Li2CT7Bv73HzXfXwAhhxXnJ2VjGtz+5QDH74V61tsyOrZ+EGqLstpwzR5UZulOcekR2VSNVK
yA2FTgi+LseJOM7+NWS7Yl8AJYdrW0Z7RsIIV++E5A9qclHfwZNO7Q7XxkJjJ1B0DAlrYtgVMieg
yO3nq0k5insWr+jpsbhcToOPwXZLtGulpvQaNNXdUnZGjhm0skGC59+LB4ZOdwYGKHsHomsFjQqo
3oj1Ju7C7GZkjBBo1FoK7ZJPndYrFKSrDU0pizqOvR3wM2/OKgiXzccsB102ZxPSzEVJdSIzSIpE
emDtkGugcEnqAi8DIirOodJU5hh+PEHwzQ9mlGD40pLG/svU2ZzOzalL02hO98Ob9HiZKSpKDdjx
4bij1wQQ+CWQz+HHm7bZt/rNPr/WeiJVE44rNgnnlC+i0V3p5SJChGKtOI4gl1wxIWxDgdNOJSoj
oro7/B9HehbmZCeB0B/7O3OGCTwIWTIUxXn6lhjPMHEJUaDscrPqflyqFK5/aMR1BA/A55a3gYKT
uQ9Gs4MHuwJGpNkaZ/URYgYbnPxUNetilW8BmcQCZxslqCuAZT9U2UbB9HGztUlHNN9krzLgM6UT
P+wptG0P6hS9i998HaYlF4ZGvI9YTqvE9CVvhMQjpEQTXoraV8G1HF0B9fQWBM1E1iIkGAqEg3bw
KRDUxn2LeeUM1wgcVBipDFogtT759tgS7DXvXdxzNRbTyxN+1eKyDpeJS6Kb8bpXf8YaZJg2UXsB
i4C177eoE1qpFscv7SX/nsxWTI+kVTPbRAY1xJcCO41xOH6c5fqKynRCDG2B0scCiK3nJ2+4R2sQ
CaICQEoWvjISzUBThmQ5KjR8+KDkbq3V2+GQSAIGYOaayaiHEulvuVC/No+C+hSuxfPucvPiXIDV
fEpNTTyee9Ec5rMtIXp374l9HlBV0UtkEqAjwLRf91vmQKW5NvOw8epYWWT7eC0W+B/VbUEnPAoA
/mTg+gEyZ5st4tsv7s/kL6Drg4fSqne1O1xtIfNNwpk9+QZRLV0wPJKDScvgWZ57HyqMJmNyMNaV
uvnmKWp8DcogyQzpDQWhHBbRNKL1JGo47lRprz/fgbV90RLU36M8f2bNH4pd5Qx+97UDDVCshGrd
lBmaeeUPyNIlHeR4iMHpI+auG8ScnHRzK04XiTCKe4B4G+Wp8z3TOsKEEkq2Cw2rmXnsDogxl9lC
d7gsh92hoaa8hvqrsQUqsCtoQkt3mUmkkou+EiorWWdcRxr/P/7nUjx0bF1ciXwe3LJB49QpapNg
WEn4gaJl8n7+8u3lRF8BFRL1wJtTMt+w0YQ7P5SnS5Iueglum1Qb2tDNgZz/AtQfTVV3iW+4fjEm
Z4I3ZThaVcCqT0x0ErXkCfhqWsPHFGX5MYJ2kWzJNGpqL+5r5Dm3K4hDwn2eJsfZsvzSGIgmHgIe
LNsSU36dJW4Ubib0xwnWhvbh0/bqhzK8zzrLifLmxA/XjzdaRZFnbYBazEZVb6QbB7ZnM/M4tIPB
zNwKr6dI6GCJvlq2v8s6unWBJn6zQ30pry37ICBsAJziPFlLX/tyDeOqc9nhpHVTUeSlGaCQQalp
qBAi0V51gQq831KOR5UUrjAnYXR3/Lwgo6TslLFNc6rUkycUwL15ImQHl1X7DyCwIYFvmSaBnZAA
GcLQFwszA9MFYy1wi69f3MrmwgTGh2fPGPidDaiXln787T009D79cNN4t3OMi9vOaCWzUaXPEJn7
IULHssLeqL9zwepv0hDA/njMK9h5trMbc0cv6UlOGjoOpPQpSxwYQlV/08bcz5U81rtwmXTgIF57
2f5bHgOgFIvH3J1wTVzxqmRie1S5gjjFZQhenoK71JSUByroSlARsQlSIf56uFYZdz25F2F0fk2h
a2z/aVp+VGOpBHpbkOddcnSyDX7nZfxqsXGWJSCweVLPkxgcgpIw4crdOMFUH7IckJTTRkB6XCP6
/v6cwSJwz2rIoG6fXHzmpOpVXH1VmOTkB5a7wy02zT5OyHhrFICK8+2Pz3XA2NYGzeWGdN8oB1ne
16zJDv/lRfthXnSRwT/nPrX2179/hIybqK4sXPNMLoHqII7tPTcmC/jZDicHIm4ujLiU1Ozg/bRz
t/9cpgGl/L2qA+/kfeG45echyZfPLuOVXw4l9jP7Sk5TkoglaIzckFzlZUbB5tP3abeT5gjyVWoL
Bkt3obJElRk4rNvl6FmolmHqWIwguKtpgeYO3hnaWh8pPE2wgLRhZuHrOa46bYN5sHhudEhthAQg
d10amreAS13HhFI6v9Eekgl1HmbRLmtfYOyUU/AypB6mTtjkbWlHq9puiryLwFaiyWdxcwSY0tLQ
ZUlCHXspwHeDl1Llh703HP/6TqW6Dop5lB9ryyToKIMrmoks/U5j1b/9bTR2JUTs1KVVdDcrazCy
S5jtLaDknBMZRjjsfFs77Ri9qLCnz8UHTiPpBIxr/0ITxzFf2aUkgEbpnPkvbG2f0RFUKdl+kKC1
YwYZ6rOc2ClN+4kDKiIwZqdvBu/fP6vpJEA+0fN+NGh+Q9ElxqzxZ/zfALDNNCHDSzCRg3K9rrp0
IJR+k7v8QQ5gS/daYV9ae0LjU0xB3VX5MfdxV8SVuMRWsT+rJNTLNMs4PwbAxtTY5GG+rwFMLFJg
hD0neLWVVolkx15/z0bQi/3FJL+NdsCtpViQs9oXVQpuc/XKlwsGRLOHj+VwoD2aw/eQrZoXqgqQ
PjYKd05HyHBJP5L93UftdrwUAq2a3qqKUpTleAVifGyxkUcHokNnTY0pw6A2QDoK88rvLgMoWSsb
mSXAAAj6atNRZ1ontTE/La4VzewCtIjNEezNDQlAdNdt7eIHX0rJxtnoAXhApfob6mqhlpEMroqr
YMPSKvQlSbL219To56cB9gaaB3B3htPpXvuHX3M67F7GWb4/cxlTqwCatMknAeXao/Fbk6aNT9nF
XL89wXcvVupQlxFq8WoLnGsQzkQrqyhVNHmXZDtWTqKySfZEra6E/7tmsqeKA+yKyRhiBEsJhgrp
jez+gYzYDzx1viGaOxSLdlWQUw8eU7V9x1PxMw9S+VlcDXzN6UreNc6qQPUKq2TyQwG4WKQP7JoH
RvpVF7bw32SyAKapNfk4kY+h57u/xgGKNt14hmmRHjRMf1eX9nD+5b8vpoRQCSpZXoM3a0AhrBVA
EwBuVhnSBJ2/jI5SJ76UHKIHIOLNb6AoU3C3yg/8x1FKNr9gQIHutAOT503lwtHdcd3dyKZpf7Ao
AmDvBVHf/a7GLAfXdgnms/12zOyaIhCVY1c8mjH8c7XWtETLN4mcLpnbvCXb35aqVl3/M3nmohHr
83qafBOun+aAB3WtSTzv4ckuUHM7bLjDdlPplB0bt8YujOKQ5tqNJ+G6/RKGZ/W8pOFKLWmpy2xI
eXH/G2cu/1fO/3x7xluxbGAIdyrR2LqUzY8EW46fJCeKGxfKZd1eLqwAxODgA0cwLpU4MTeUJz7O
q9jrz3AtGmo7x+vKukki08Lt100RTiRKSsa1yOSWHJtxcc4YvYFzX45fHOpOL6xZG0nvhN9tIqF0
3nNU3mNn/kwNWgSTcARFeuFYMv+eo0CKKIozvIQtcU/5pr81LVxmSUwqtt0hu2KiynxucFG2DuW3
N5O984nKQdswD0xsBfkwoXBh5PB8PTGtgA/cfWyWsTY/IA6vTtkB6eXHkdhyZTYbIHdnU04yDcZa
UslrOT1XMVZ05ZpnmRxskwlh0Q+MndiR6OF4bDmRiJvKqt0YbEQlDnqtKW7pbwHMeO3ouHunX+hW
sMh6xkb4gNctPK6GUgxVQG6sbU3sEzxYUTBuBTxhYWmUrX/U7kqKxtPirxmUO5+S9GItbLYaRtsd
MqJdDaCWG1QhXSoZ+vY5hAgwXImghY994ZSoD5dmP3NIDl+Zum743yg9gvMtH3fwuFKSIErNMv09
YePswMvU36J4zqiAK5ahm8RJ61M1Z52pcHhSi+ta2L97P/9iVjtPmg1pxG0UntbhPXGO6QaiizL/
5EK4DWQW/+kfxAmPV3MiAi/f6KuInhkvi4cwJvZadnJBVWOVALmnN3b8Jt02q3qZCPdd7qYtpBcT
gQNupGuHsGg2Jo5vdbWSyN+c+RN6TucwHTwjLROa0bvAC6SlsVtyDWxMmdMBT2hlX/XiLqGqtISZ
Fe0eKH1jVaXSlexKaak6l9Fz8o0DHuwwSEtcIkBm2jKKSHjqd1peXPtmwIODD8sd9b3mIGIDHNDA
Sgi4R7P+6yLSkI/GEA6gZC2JwULg8VRp6spFA1mBj25KmpBrx3jftODGoB7HSieaunH3wxcsLD77
vAh0OWmQUS66tXyzs97sPX737pUkpLAyEBJ6ggZCu4I4EjMYrWPBpvtfsxmiNyF/nvlvnXj/23t2
EXxpyJbEo5CC8hdUPlUXzrSXPqggjXS9Qoha8wBCQlpqLAVEti5MqbYnw8l8Fq3+0KJ5h7/84Tff
xi+EndUPjPLQ7jPar6u537SYT2RSgFT3u1KkZQ4hFKy3GgW2huagzn90P6qAov7XIt+UYV4oy6fa
bnz/SVHpp80UjUGI/oJgDIwHXp1c0qIj5wNTwo6+8XhVf8yuVn127vvKt+RyFCra11WjJDKbqBhQ
5TLHRL6oBT+YxZ2Z5/8U0NAasJ+2dPBWR+MIpQSmHC/i0XhKCwRsErGFPRAx5hKpblGeOmPzSTkx
+2sitwFlBoSWuhv3Q2pKGBjMjc6nCyBqis8K3SKa+472kWJC1J+bCwvuGmaONlTmssGkLBkTdSnU
rvbkBoq+qDFTj3yAjd7AsE/it1pMxRUvMM8DIyMT/fawpnSjz7Lfk+jNsfHZKFmYIYkxUMaoO3Cz
HIm/3qctl3ewoe7WxIxS1AFvn7d/0sAwkn5Lk2gua7skWvfAQjXMAl7fuHwyk30PYDwLw6SaqN0R
A/agW24Z6mHGh6log6OrhV1YMncbz4zhE48QjQFolvJfVL+muuZnlIFzWk4GdNO4ZGWsx57W/oRW
ZohRBmP2n9uYzJDeQFjNhq2/a25iWoTYhz2a5AHVThcSDfiTJGq/HfHb4nmPc48cnSj9aCJzW79p
ETGHEMHP+zV8PZ+vHMBnOGm/XbiDnQy39yN2k9AF81G5m98Q0xf+19wCdzrOHMfLFmVI24U43aZF
s/NHbpH9qzZsqj5i75tCnrPXxYEW2ItRprkRbFIsyv96J5tximdJ3RkSufP9mHJV25QO9VgOTfda
A7JU6OWAlYftNhs6OIt2dlar4DyumMd5eP+A/GlXGLBLxt6JEYJERpfwvEBeuCMRs1a2YHSxcdD5
05KCjAiZ3H6GPF8+XgCWlgG10ZEZNXeHb2kchQjzRa97t5nujI7gtYZLg3zhcTzEIW4rF0kiBWUi
Snn6ec694TOvrng0/+NcaffoBLKM4Ed7jxhwn4MhaWAm4T6MN4wCurj1GR8Bp7O1JpPV5Eb8hipI
hx45rPZPOqA5IUKWHEyYcIEMz/nqgT6ftHaF7j9EOEn5prX3guIVO8suEQRzZqEn/ms0swyiDwTb
GTpl00FUzTM2eYl+uCh/B7Mm7x0yb2/X/Yol0/Dg873FYNMZhEpaU8aNJVk60J9HS6fKvzEkI/6e
GSA/amtqY08gNlLVbXQEZXu5CIDGeTuH4NSbNfc+ZGq0duhYNnJHjmEfNrlcDG8wb9NoV9YzBtIj
AHBPJWeywzgD9DmFGWcdqOcLBXWqe7rMzs6PIjMQa1oyETNuNrfUDDjDnqQU6rY5Z7D6DxhVfjvH
bptswRqETB1s1/nEFnZEvlcs0VhenEAEpmR1aV1gI51G9uMz65eRm1fIAu4G02sFWjXceZOst7BP
AbaxlY5Mb35YIAsXfG0VWHdJvpBgfRCtOsE89VMGyFdAAbl8vzvmPr01JjINEaN6RoO6JR6572p/
reGdwM6FmIAbuSiJymT2a4wth5RdJkvK5hgAjTBzkIdaPxMqYJiZFuMvhV7WIyKtWdwHjH3vZb+u
YD9KZGoYSj/oqiPrW2s5I+bEwtvgfHt4iGS07IygS10kugya56DTQkkReyCYnrXw6xdiIvuO53mS
KTjzH1WbEw+AB15n4PCiYy/72/Ump7g6W05vhVvn7BgF/AvGKh7NeZRk2BYaceo0IRk6ZbP3Vcay
1a+26NqY7f3366I/0x1xMkBC+AcvcF5yHBNhs64mzV5jpQhdTtE93Yukmj1tgNAsmvyqHA/w6rvK
r3+aOIoMQIVx4BZ5BB3e9+DYcF9IXG7/n1MKcblNWjKt022bpD+7YPjUM7l8PWPFd7q/rq2xR9nm
qBtJrDz0Cu8ejrk+V6hC9V0Lb/tjdHOTfOEZHBh8RsvO1lKLwqO50t7Cx9pJj6QjgVU2fNveV+Wc
diWBCGhfNqStiygeBqlvVwssiPw/zRCI5FyxvbFNPoAodRnejAgd7Ax6NidyMTZM6qlCMoxuCoZt
GHXVuD8ZR5VZyWXd5BGng/+OUPOc7P2fVDBq5DemGkA5lmwDGm2p+2DQji9p1c4oM5PQPXj6ewaC
R0U+dkmFgoMpiGf6DJ8jGKwwibQsLKBpzhLR1KHrtplyJkWPoOlKSUZecbFAmp+G2GsavQKGqpJ6
RDKxVY48FTQeo+CsajU/bXanEmNZNzuPiKGv1snnZxtVo+LGR/k+kKLEgZAYDpFfpLrpKRE4RAgk
4LftEjNMfyK1EPxVUpV8DsZXRoD8LK7YLxggstcBdbvWi6VR4mksaPZDxholEpW7A2HwyaPRE9Ti
dzVLxRzl4dE4L9cO1U9JPde7ShIW8ougPxLooVfXHbr+LbqLv77KfdjzXbArYCvmEhqQh9UVmXpi
9K3IGkhvVO8r6TwSmUfuplXxT1rKZLIYxGB7lc4ZsYQyYFw88u62UN/8mD6oo3Q5FYeibTU1tAby
yPfSqAAfRCNEFVGBta54wsQvYqbrphXD5T5RPXOvmJSrqI56FSPYcoC9FrwpebFrsAjqNMe11Rk7
73sH+RDhcJutxoY7X75LC9DoMoxKZQyJ7Fh0RqoaKeKyY6fpKu3NID6XbUiIlqh8K+XPftDKL1KL
gWFVqDJnNjSDyWlwFTMiqs6Ut7vui6xmNlv1qI6hZVNCqZu5dvZ3n5EKXPOVMFI/Gthyf1aEDaa1
gFiRdovXNp0zjXcarefWueqX9tJsaFvYN+C2pPWxZZXLdJSQctZdjf640waQa2/vEmwrWq3ESliZ
H7qbUlBdnRcO1KM2HTu/fb+ysPkpq0L10ftXN26w+zCj+MmCbvE+C54oSf3Eb5Nyy3CqXiZl7/1r
pRDTU1NMo5C2XzT/6UNKPNbp62DO0nWoPeplqPdrN9vAuGG4eQR2iOLaa2PKYrVzfqZxP5epOrnt
4jIi6G5uNnVrZ8drvZrjUf6p+ik5Xz9CQJUU+2agC9lGOzyNSkdEf0dq49Fq103nDfUxyNteUkCt
kTLP7OtiCN+6NKxjwzcUIoNUUYGvy7IIBN5fFTvroMODBSM19/zfZJUhrWlEjU4TPiHbYMCu2ztM
quKdAQfJJ4InbfZd8w9pJmPzEBiXSy64DJUWRUqiPMaDFRLIauYlh/vUbjfxu6TV0eRebTbCd3S3
TlTCiF7q1B6k4JLJKg5DoEtGNT9DyWAPzQdzM5RKGAOmfpZ55cgs61xYF1B1zyI4VU0x2G2WIRGS
LT0jGgZRwJEO4GEl+jZqguUdjSErQX6Jtjlz0pntYI32/6aHzcN8vkjmCT5tHrT5n7+SqPD2f+DL
E5ubbUZ/bPeOT831LaT3wp9hmkW3Pf7ShsXdFnHgPOnzq2puEBxc3lqZ+PD4UhzfsvP1vuSQktlk
r2HRRGKyaQBU7/dwUjLY5LaaWcg4u0fVvzAD5zFA0v2LHaqfzrtK82f1g8gUfDcm4nGV22qQRCGX
V6ljFyo0IvNZsXcQ95eyf170u/kFw+VvcVT1jx7S9L1TMLf/cYf0mxD0ko3eP9uI66Okf6qIAijV
Ws9LQMQ6eALx4s9Vh8oko4+kAltmc8bxDTqP8eeeKNwLHsGZJQKwElhx8x+MWwnk0kmA7NTaEu8G
vcX+R0Ic/3Q+Mpt2I1EsWDWDIDb3Gu4U8N0mFW/KjixRY0pMz7AJQx0q9mSaiCGiNsfGLxaodDfA
TOBzUkg4xfwrxV8evRQMdd+Iyg1jQbnO1iEV5oWtcJsg+pjA4r9vuM7tmn5ClkC1BqyT0gJUUzsH
gPsgpuaMBR0Uu8ZwiMjKnqkKFHjq9BQ12PaHKVmofYTG3OEwDLwjnPX39Om5QcM8C6/36ulfZy6V
qQc+s0tbbay2ID5txOxbb7qsbS4PcKxe6ZZ+ddzH/wh/G0HPTDzJ2tlxg5vInyQ+6OK0n8YONXZ/
8UOH9eQiFYz2hN+lpEtG9PN7gkMCeiteVJ6ZopJb+nMANodk7czbeu6t31YMzWGLFJFfkSMWttjy
D3C0+y2QPMHtsTbOx8LChu3utYw+GlyJ/NUTqlfvGQ1aZJjWJxN5WtEBnhf9OpQdbmMsPRE8LUFA
wxnALmooAcV0zyTae32aZzRfKaHLhBv8nHbFF8MCKxwqr9A3gkc8UcHPJQqeIBSbLpydXBQ4eJb8
ZfBhJ0ME78LRJuXDNPVk29r4n9pxjCHU2LHl0My1+3LypSbjniPpMRdSxEk8hiajWkjwkaWS4NS0
fYKw41r52yVPK8AOQeheVuJDQe/Ubx7VcieT1xBU/2QHzy10kwF7Br2Buj7FM2h3L2+MLAhotCYf
gg6rIoAfbpBNPVJvbPgu6K1CYTYVoIMyEmOsfhAOU8vj5Rz5+821BP27Q5E/A1on4X2QtHDeA0iE
wj9a2nm4UYgfWN08SJsFnVhmgUn7LXwdz9m+HjeZzX5mChlXB4n2vWU+u2FjC6AxbwjNg+KXKQdR
wUsABnTbN+jtAk5dpqeJfPjqb/TH7EAl6VXpLTHH8fNgRdtoi2qAYIiybf+Hc75GyokuuhoQwI4r
Zf4i9uLoVo8C3Dm1RmdGtL+PmgB4oeRADEp1XX6BqSCvBJ3afHi4LeWjLqqBzgdkxHBBCjtrBBru
iEv89ro8tzR7K8i1nn84BQ3rCGsYcQXOYO0w2lMKAkYAO9JsyPX6ZHkxfX2xf9I8tlkfhlAQCKuc
LxoC+fOHMWNxe4M6NvDcEEf1qfHl6DwEBWUeVAONkpuwCPfxcfPsOsdX4gzKQ/x1YQFRTOO63qvl
L07W4ykTziZAAZRux80RJYqRZ2vAXk4GYh4iLEgzozYprhdy0Key7l2IlMf1jNzWDFSSbQrZc8sJ
icoVqSr4gZHA/YazhD5CY6vfoj39wHV3pptJsRw5ctsdXK1V13UeOowNk1cYnai2ttQ1g7oW2RKr
QOSx2KRj8B5JS6WfP/HCrNiMRsIX2zluX4z4XZI9tJsM3Uz42WSEsPol9jrdngIdlKdin6SE/HC+
CTAaRHvuWDtkNvsFHiyFmM/5KoMQX6k0QQRjNdVZ7X68dcS3osV+tUrMyP6ulgTWkc2Z72tAj7d4
FroDw7OJIX5wc3guiHzz/ULJIkqzWZ76dFImkIu6P1jU5FVICiXnXbXoTgShbZ7YBAs7f+PUPp6K
mSDpHOPwGmWSUhSOdC8fYocHYIN/LenpBQkexU0b4icoWJn2fHQEHeNsjP0Y1uieyqCoXtKWAJYd
DZf1wlNiHtv7qMoL2ssCRSbtmTvI5bgpufR9mF/+R6v/YdQTPJ578B468TE47bcQ7sVQcUFWxevw
jlIdp/j6F4P0GVrbaj4OyUfn0ZkH8QvFCvIRKJMFEc2yLH91Rjme4ke1Uze6NkZWL2+o48RcdZRX
Xk+nUJWuglssZPvVDJfgZDZJJNLtpvgvRFiQAz5nXuvDIH4h7QJoRgrGi4H3az1MfYgr+n4t875+
e0dDxgW3/TS/JeuPNYxshtnTpaToDRA1Fyj6xsMtLwFkpPt5M6Y8qwB8+6DQe0Xvftkj3NW69E3H
RB3A5FcbJH/CDn/7MKSXnR2YcXqtDxffB82IZL7XuvoI0qAe7bLKOmGqKWnQiOQfl1MwHctD/W+w
DAz4uemTZ9Fn/hZth71Av08XDJH+0ms+N7L7bBfjt6do+sMdPk5Qq762VbdR0p7mU3GBsNQ9MXR1
3FxGWy4GsEtI8LDItOz63AOcUFgS1RrMS1M9UuuUtub+YEinLkJjpsd8JZzMUA/ksYVjugPUBM42
FclfJ3v/Mi3adknzbUvg4pxjC8ISjDxereFc/YmHxu4SyqGdouxMLtNBiQLRivcFCvr6EGna0XUJ
y0y86Ld02VN5QbiwX6qyZ6IP+pfXr8vCf5ACnoGHxb53aX/ubD7qLjtFACb6MZPEnDDfecgV97G6
o4l3yJJ+kAnzDqoGxSmnyuTN25pOjKGBZKhdN7lqgCAtBIFjaZ0NalI5+19Hn31tyWGABgtqwAj7
QnFjgmW7LyhhGqFedzVtOZfbxv7osNsuUzEC8UjdZeEOPoL3FJzt5VS7vvWtF7aeVK4XaIlbe/ue
S4xrsjWTaFcowmh3b6sSPDql5aoOCOrhZ0ZaFySTilkR+5iihi8NjJm73FXNn+VkgkFQaIAV6xWh
5FojPgfEYmOABNEKEck35/bN/gHU1qPt5W8mu/qjBlGm77B3djADHt27SmrdsHqsnH176TdQlQD/
JX2VPJIImGh0A63DzX2L522F6rtDzJx+bndriL1ITbE4cNFKVAUJo6m6guVj9ljgvtUjmEnDmOyC
Ju9KOjF1y7dwSqid669tMe2LnoB5hRTxBKDWA7AcZoDP/Yhj81iocjGfEYQWJGFJAMWbDZMTigCF
cCBz/oI5jV5/o1g93fm5o7Aer0thgJTzIJjwTGVFbMBtFPjecCNR8ojsR+v/5WTIrB6YmSb90+OI
JJFH4yQZmtMHIIvQomF44pv8MNeAhtbwKNiFTPSjfgD5Jiwxb8HROEIrMYPlVtoM1Ezq9S3IkeYP
aZOKzhdq0LVBnmAhf/O5+eoCE3Ue9kc24WJhWYCnF1OPJFDcgxudRZ6Iav1xmyRcu/OSvYKTz+j9
uJwYVo5pQQvQBJ33xGQxhUVIiiRV8DJrLRtl1S8bay7oNYrXg4KoVJgzZ63NMbViAuykkDnmGFMO
UHDXUyNioRfa76diZfOExdgN2Wzo3O7D/sBYVaMEJ7btbFFLp/bkm4NXMI+LjoXZy/UmbywUIsDi
+gTHcH26qif9mhOKil/ZQydueR3igCSAGgPvvHrPznxQQmkXqcRGNClSKcBVDJofAb2AGW0S0v8u
vo+NmsNzipCE8p4tNWA7qTarbwJBAp2R8oJE5vKpHMahdUgpPBM8xbZVgdlpfvft9JB7rJYeJn5z
G4IASjaN2/o2GrSwVLrEwQrTwPPCeqF4UI1DM+YJ38dgi5J1LpP6l+KwacVLKGxGplYdd5IX36Jt
Xf635yHkS4+4PDrh8HhfQNB+9MwU9dxQE0acQmkt70CBioR7GY4byEJUfBO2+B5jWSNUl3Y7Dk4k
Chet53VX2AFOreCHVr0VEzRPZuQb/bwhbhVr/L+4ZudIL4/9S/70sDs2gfPrt+y1bT6QCAc9M1PA
A10xKit0ioikrYu5SvGYdqM98lJJiVGx4P/7YkXy4krTkoBMeGsiMuDyMJ9VDABXWBZJXQDTXooR
30rurZUuspfvqaeVehh0to/tp29IcwDOWYGfDB3rml3IaFEaQY3hCYmUnL2BYFM4jUPUWePNaexS
k4MxYSYkVuyUE9qxft+wQjW/1Y1SdIw/8WZ0lll6tHwvjxk7mUYWxhlWhAiWJiO+YRNyVvJxIEVU
mdU+YXlom7nDeGgXoQwKw1nsuiKoTG3FzRLm7cqg8olUnD/L7lK1hbzfkTdtmH7hq5yV/Iet6Rwg
ItDfQPC+O5idoFi4/Ef3NAqj1buv12YmvaEF1blq15dfRY3l0anton328suVSih0mM2nTNdWSXxb
K6qdp59p8+OvK1lKm0vPad2rWK1tSGot6PxxskJXc0I10JRzOfqKZSK5o6f3W+xlPffNXNkpq+KJ
gVbHYEja0oJdZmn6m0I+sv7iL5bUcvo7thM4QHoFpjbQJvJRgtWCLNyGLFoBxj3984kYjf9xyK9C
SuzmckUsIaQMarxHKd5BBaNGAhNNYNsDx08oOwtNEMqrIy4ZTRa/QPMhXdQEm9n/WDmn+D+eVe0G
GhvKLPIXlW16BYVaF1X4uQ/t3PAtQ6KIRo2LewPZQrAlr3fdBxjWn0C+KenNOiyc+XdgAOtykprG
tufGSwNd6dIPrB/Tfh/Kt/q1NwAq91LRmsdMJ6ZCD6bfWJWWW/tRkUJQ7+5iZBg6s8gdglT0NVHL
Y2C9SrSUKj7GlJ0q3tg2rI8ejUG44Yy6V+p2zAL3Vi6XZCFjs2O6YeBGaCp1JuzTpeb1qF45UJqU
gmyDJz/o8wJDRAjyUYYTPCAudYz0c5MNumMGnaPhOur2n1aYgSKqM6hJKhlmIyiDLfheKcuez94l
PrElYIXCDn5QL0RbHJ+llfLU+T3rGNmQRMQMK4ocTGQI5MSoU2tEfMReRRJkdbg+v1Hz96c811ND
ceUoY55ssw4SpisomkPZHVasUrNxko171cBnwi6p65sPdH5C7JFEoqnWDbNiHanKFJuW/fN+5IOp
0itxQlWt9tOzFlrvc8MbTIv+Ac40UHPdRbfyiqE7DtbE2c+cSzCo809x/2a7SJSoFhnZXSDUivmk
u15eowOlkYtCBSjdxX8hW3BbnOCLIhbktnzejGkJoSh4y5HWitFyGtW5/kv4XxtQdZyLth0brIUu
ojtRbsV+z7WMtfVZ9y5BituSHbreRbjop4GSiiCHHMei1SELJzFde70GPyyB+bDet77cc7M1EhsG
RfXB63aIfQqZT0iJ+BkcFodWdOqsqgmirolHKi+N0PfHRydLA88W82x/E2zd1mEYPEu0cvn2C7K3
atoIzfriOw+ZMl+eCLCjsTu7AoCuyMgRqFmCMUnVWhNsGK3B7g/M3WzEd8ECw/pRQ3D7a+3kHDqh
lX49PIw2g7JaLLxF0Zosw/hiPgEf2vvdRUOdyzm9xhxfjVZtOPv7eDHlotpLKhTIPPTkU1RBU2Io
ZXK7vrVBV8IgMEx8E6a+GJcFGl8JMr/NmiQ0cfXxv6PloTXByQEujqzu29fnZQXLOCcxDPxLJH/j
Sk8MuCI46kzuZwZ4e21qne4yZ9Su91Rfe5pKbK+JHsKuL0sPyVZ+dmj57/LvpeXHMnbqAVp6aZtZ
FF5UhE4fI1mRh86BUE7El3HUXL4LSqx4khqVwA10/DdzuzAJ7MSdAZud0LBU0yOiDJAHVQUNlzHL
Dk5MEFiBSb/QcBfwUq8LgyDvBjwULKGfGtIeqbOHLEDH6USGXvtcWBeZ/KT3kcEb/pwexReHVY8L
7vGMLfNW/pLvrBVDIDhuS4AganJ6u1TUigQcRVAM7gF0oS0Yxu2MMl6uNiJ3xJUZZejFmKkGF/gy
76SKNAGZ0P0+r2XJm0OEQBEmZRr1ojaIfDgnirI/vCuY/ekxz0ALtQoGly0rn/wLQaiwFqpbzg7l
2XJOBCRX9WCDFmLcnkXR8R1futhTKctj3duZGiTHOr5Ir3wGOh6unOamnB0Qnxkykl1ddQKBApAU
U8tGjHtzq8b/QsX0FQQvht4eOlYxEbgMasCN2HiyhA4YQhg0GFdLUHcRGAzG8J1p+UM2DYjBnx3i
9K0ByejxJbDRYp8uFGuTpeS61LMlc+jgLrj1LCuK2GgjlrXPucSBTwmTaAp2lsMzU0+ZT0lXXdy4
q4bPi5/p4IVcIexRFOaz5rCGwyZZW/rI2fa6cbvb89qIvbEpoU2l48l/a0M0ge/LXJhWMgUf9KzH
OS/VL9D5l1S3RY9aDx5Uz9cilVB1Opoi4qh5PABKjZ+H+acTwYa9QY5uFVMuDCr231D8V6eXSeiK
Cm/JjbhVs1rsJuCDbbuGRzJQnSoHSCII5rA7gpRuGNcXyqVKvL22Bzek+U0slVwz8iRoMmWfhMjp
IaV2/bmrn4kxn+Rs17ICKAhHWYpBA5Fu0+vm70dlBolvYfbA/gnfIKswK+xv7nF4wm9B1rNTnP9p
v2T+iYcnsVpoQN2B7X0FzAi+wqmLRgfiZpaRcXF198CxpZbbBlGjv4J2tmgzdwGVuRnlQTTb1hkK
jYv/mmxCT2J7WzOwWQvE6SxGfuaG4Su4WuPrTsMEVONxzaKTiqOKkYJ2hxOX15xRuI4Lsv8oRE0K
2e0KO86RNYNukavx1RVDAhuN+OZ7iV3EnAh8iLv1max4uzIzkWI2Sn9cxM2+rmMcpl0o3e8ISvvm
IgsGOmpFBbgS3eKkigB+sGHVDED3CQg552iLJxWUX2BzqAnbBsLhMBxdFCVkFTFPTn/1mVZ9m9LA
3/ckOBpk70BZVqL5VVNROhGswP3M8G2qJNE589ccd1EkOaxjGvLzKNrB4o3Y4pHOeXScCnOTA6Rq
Grs8WHMM/NP6sM8UQggquhmSvAhwgq4s9o4X4dLRzCsl0OApYEFGhRgxG/mawt84q93qoHRmUth7
Y+BHg0NIZfuMwE9Eq55/LW1ShJklcF1U676HLlMX+0H1vmzzb4taJwpiYB6uOvnaP/vHdHpfUTwp
qJ85rD4MUARAW11OGdtuh3TTkHaudp8LB/FIO6wDoQVcwDGnHQKisKTUoWj2SIqbnDrQiUqtcWQk
9cguITVj7glmEYJLI/90Ce2ntRtcu0d6rpkDZ7HkkYV5sRY3GwCNzUE16eDj5bLjHIBFUTJJUflE
aNs38mCZMxAgef9DfkSIdGq+sJS2+baaeNrQ0/7i0RDLk5HvKsyZSwxUJcvbMUf/glswMSH/lZ9b
8tT8R6HSmuO0agpg7YWjxO/wtqO4efSH6xVgDrf3vHxiOxMgPTcj1ZGMtrfMR2Os9IdVx3vAG3hm
XuW6gVLiCBYs80ZmBppsANkZTS8vgag4WqfrLoVlB14jkK9psFNyZbJEKhBd+UCa7VtUapkHJ/LO
6zfSCPEWOZ4eHHa4G1jnVVBK1q5P1/lJNUsa7X3jP5cwXKp/6u9OzzPxO/13r0Nf7XfjpLM0xYLp
fxj2ljZaipUP5MmWRt7nMfdR8B0GBHTdNVNJdpn8s+/W9KSJe6m20kG2rI/Ba+IBkmiFpGGAhpIo
og2+ZJ47HAkiyPIfX35wqt4fS7knHj3wtwhJaWvarJzNDtJ1vreGN+LoGdqH8z6Hx0SMJJOa2dlW
/ZApi3z7Z+054y9D5tz3spc5hBkTaBnTJAvu0Nz8646q6Ut8UElsNgbUGBMJEpQ92zgwd20C4NuR
Goybh0gC8cpvJYLiyI6/EfyfdTH7OIOGGuKmy/Wmiia9r55ge9Nh6kphwVJWxYurjDwVn3objMFA
A301a7U/lMDbG7/304++2dW2F7V52Q48Yu2Pw+rsCFqoK+S5gLk4u8BaMmgRjlMJEfu0tmiztZBf
PN8pO6U16C+nhVytCXko9Ea30kYlVkYgzRlvHL4+FayIk3LIHmFeJ67aY+Hy0jRuhdUGIEBn3fSc
W8inwDDdPyKq3DaQFb4LBQcfZbqq6oCupNp+LuHNT0SfCdT4JM87l49lCLLlLEC8JPODN+ExGfN2
IjxDk+AQ1NlJBfWMCv/V4P1TQfv+TyVGIiiEckO3ZQLNeNS/n7lKJjcScxkoOMB5CMrfqQl8aUh5
HqK5iJivU2Ow6YoOXXDpzHnMpaiorXxxzMGDXXHK8svWb3YIYJ79hrRbqdnQo8LAgOObviU5F9P0
UzivEgGtwzaYmJmkYnM8ZsyCzYS297ftnTYCsEEubC4YFFfkx05Wg3BNRDmeRjrtpHnznoT2IeIs
xxiX3u497ZAD3JJXUhpklf9XirrCOqA07Wyxe5BoaQUWKKYM8LEo7ZgroiCjLzL9HQZG90ntd4FP
V8aU8UXQrkVM9OHYyotBu13ToOMogcjUatfw2Qx0sVUqWF7kaWyv0qr6p41tiCfdYGdijiNZ9WDQ
q7Zx08+2ZWWsH2ibltLCcViQNqEVfEvyy2wXdRjv606nVUqX17hRYxTLzjIoUUXTQlFDbG+DuELu
e81VvJA4nIMN3mU9WW4Yam/v5m6vGZhG4jw4LxVN9WKzT1J/MOeIXlObkUj/n8wwrpu7VybEdOAW
FNDeYgYwZsRIudVjYoKaTJW/Uc4wyQxsev+J3kvonRNXemF/JB+/zwuX4ZT14XSdRrvZUdYsPMvm
H4i78vUv+RyeSlvqHYs9tkguKyq2Sh10UYjOHukv0/sxbwOi9Rezx8UMMc5M4riTYmfw85skAU8H
vk/u6bWUSTQSuusV3rL1s83I1qACkaiXGq85gdSqn8OsXUM1AnGRv7WFSVK+bdAwRMvwZHsQ4ltT
4Ve0D63EUq/qVp9YuMjcOMTk1LSkcxZmQwxMtNuv+DR4AUGJEWlCGLjIMqQd6D0plLeZl6PJaphn
V1dkUGZ8aFIhUlLTcVT0LxE2yE6RhmSJTh0G6PXQxi29YIlTrm73HOrAv0y0uUixuzzRoTtaIjJi
ok8+DYhHskK5gPSr/9HNhJ9l86R7nUb1bIdt9KfxG45XVKnY+EcpYRxF68Z8ZXCKD1iayD8CIjg6
B1Yn0N5meYhtaAuLI9dpm1R/B7fwW4UB+YY5r0Ef00FnOjyjEcWi6IrYJZq1bwK29/+FCe09+37G
aLSrqJZ7HUhTZJ/s9gxUNqtMLa0lp2ddj9xa3W4xNeZWHilE86XDWLpUTZAZIpLlD4c3QqeIYlrK
+UrspiwcJXZg4XlfIhhQhwcRlMR2pCJgsrpw+W/bIj5bnC2/HaEgPQd2zEkKiuV2NrSOpVIWrmC9
ezMSnY1EslnH75JD7ER/GcqH1AGmYgifu2pW6ZzzHqDW4OhQVJTxydc56xqdnygdtC904CYxEkJA
b6GViE/duNoTbq3MGEXj5cT5zntPZOPvUYNtcR/tzK2fMxNMG29s5QQWyy8oHBk/V8CF7bRi86Gd
W4+LruYT26QtTpgOZF6mgvJwnhxvm1qX0Oykyd8wAz1pDDqD+IzMNG67VNU9agbtUndDxH2XJ+Rm
7Ovtg8gMgPu82OatkyEMJaSRfICo6EEFSgYK+b/xkRSmrIuth/0yXwxVr2wryDZeMSXpCiNATXgR
y2n+oQcKFooVuknZAVxnN478CN8mkDT5WD87uNlPLbNKNUsr1HJM8tRabjhDJsDPOdh1dnRncZ5I
PILuwDuaboMT1Yiwo+ZKS3igHoD+06myc87EbKfNQBbLtoz3+KLMlvA72BPD3kIeaNhBy3QQIRcV
q37J/sDJ2TnzvEJ2ddmiGcc/W8gN/PnW5Cdu48oOmLqnHqpxNVNJVVZdnYOnXC1i2/yUd+GBEvfw
zJGK003x+vvdix+9njii0B1eG7GswnpSM4Pi4RyvN4hP9nbr7H4dkiuu14ksQuycltGvLOeGeiN/
+vq74WvJzk3qUah1veINoniY+jQKVzEayD9oKNZid1k/NfiWVG6fYveHU7NadzU7Qf/A2TSfhw3d
2yU9mLnE4l6lkFCtyZj2lF8EEo+qZ/b9uo3GF5K7GL/GkHfUimcMxS6IfPGparc2gf2V1v7SmqH/
G71OOf3Vr+hbBBmLwLlShJJcww+GJuj3X7dSz4/jysAmsbaAsdfqJrXeFBK9rRUHs+Nmhp2mKu2U
/hnw95ObHyKf547KO2CbCxV7jTS6C+Hc4Jz+KAp5/vYLy17xeAUCe2cVEEGkHSuuSKNN3gH99kwC
TqBcVxc/6AN6xTTQEkuRtgVYWRjXMmPS73TWHS4G+aWrpBy1fWfxxzl2Jgdd8w9MfavqWx9Pa+MN
fN2TyA77im7OwSW4AedOyfUS59STpsXIdYe6/TgEbv5QyrzLpToA77viBQdOBBAzapm269ZVvxC8
xjVv/T0tIZ32SAf/vh2c90tfyAxkK55Sl/IcNxpJcdKcmOMFgW4Ojg3ygZAesZLvXAvs+ScMnmjC
1Jz9CqojIsb6+Lcdm71+AgD01XppyZwaG7XwQrkALe7ByDA5S7iTuOjs3CzZBYdzLTGW9PVdmT8U
FGnvlBbOuxGQwWzi3VM19UjvtoPX4fBYMRNMiVVJc5OAaWN0CDIXLTSoIbYyQz1oDPG8TSPyz4za
sZpw1jt/dQa7aX1Tl9aaEOw0guIY6zir3nAs19fW+MJt7djvk8/GOhMSOfWeAmIuD1c2QS7/KOl+
hfxk+4FfMQtbZDQEy/1MyEi1r7ctgW3tyZTDCIPFVCVk/Oqqw8DnvLZ/+gWTQz2gdcKmu1KIxe8g
I4fQ8NX9zvWvnS8+40DqBxUcAVyvLasY6kG7dRA2ZbExom/ehRh3LsD0smx5du73PCOjwcViFe6h
Afc/sCO3EkGAbF8xlCU7JT42NJGO2HErGV0QtqUX9WERrPypyGfUf6ZzW71T5sInc34Cwu7JWYXe
7kT8LqEI9zaLbF5j4La5K9hQGdzp4ZPLaLPh4poxUcggLbWUvfqpA6XMpuk63UBf8sgc3IqaVMSX
TXABT68mFbBoonu88C9ghofJhG4Qm6n7MR/h4kHKb1EZdA0TlM12AXjrFRths0gO1zss5PIgP4l+
SIm8OW63KFBAyoC3tPhUdISYwpJCX493coYha+vajhptXeOQ8IqltQg9L9VjQKK0JKKxPFJANHR1
QApuLD5FlsQq1501CvJfDzdT+HKcn6Q6LyRf8u1U8/KxU94OeC7AYLvmaY86/paHtS+/c4UshGtn
bICGLFk/9sRVriAmim5I0ZRBVViwRZ9ndYpeUAkrKWO0bGJqcxUsiWFzOZ38OnkBXlQdGREGT3yl
jf6y152/gwAJil6djG9rP2rdk3Zn69WEJTtbfNtlA5JJe3eio/mZd20ZjGFlt8F/diLOszXH8MpE
iUUDYFTTssLEhSEBFobmOSixJ9nGk8NGjpB9ThpwCDfnemzcM0XnI/lXSaOHirumY6KUDuUMom9i
pcyo3HbFfqiHii3J2wfv8cM5hbQbgesR2DdkS74z+Ak7o8rH2gtfj2yz0VdH2nWp8A8In8pAAcBo
yP9i9biPfb+e8RuASqzP3F0Bl0e+LqfzaH0/au9/49TPWYZQBL5GFDWt4cpRSa08HXVUdjZm7Ch3
3CRC9dL6kwk5cdm2A22sW2kquwLwEYwn3uwK9ZZdl6WCe7xsEAYcgcF9rsHrfV13597VM7azSb1w
0ICbcoMNM+cx64k6TJDHxqS2K5zIPVnc4r5ZLeRSnMG/jeW/e0RrEyFevkUXVqg60jpc4zfAz7Km
fK2DZyECT5DWfPAGR+HFRVvsXkTrTQGkXMSvZv6AoGdg0eN1CoSNNoO7FF3DyBn/E0E5dijrpC2R
LhsZA/fBzDpT/y2G7V4sdxlqaCHacniWlKPAhdvCpn+gKJFZSp4iZ/sZxXXGQBvY7ucNAIDUStZQ
iq8r2c8riwupXzgdGZXELkO81Immtgdi2Md1Cpn+YokJJspd2ZSTRhuJaFPI9H0WTXoY36myF4Jw
XI+6Z4ozusLeEMb5jb706huB/hwtHaa9GrEfzv769nsSM+vkcy0ewF+PPdvaZIjnZHNT2VxFXpDQ
uk8L8CHMnlRrMwmsUbh+K6xREVGFsSYLoGet1g8YMdgm8VHiAxFsT5KH+AI7aJYiCFbKxT2eHMBD
uQlqbF9cDddXEDleZhPQxGP1roImQ0Q2Rp51v0oKwXgsoTpyvjIvaoBWzQPxfmUYICbXlMWyzGUt
7kXpnt34vk2Jop+aQNpfL+CBQXS8UOJ44I9xoUx9MYjaxFklHLF7QSj1oi/hD4ai6gwAdcx3a45c
4H0rcqAfMVYsykOywUPFTT/msXh2L0GE3XRUhc37asevCl+AhFYkcrsig/iuh/YNWK4Dud39jGh/
oDtVmpBELn1vGXQHX0aD7PUfSEdu6rTOaZCFdNVt9OQ2ItNFowFDyWLw3dIVZsQUOv45UzIOWLF/
a+/xHpWie91lR+f7mw8n47Ob7VFDS+40PVW7eG4MtxY7+Ceglfp7LsuwVOlBWTlpWAI2EDxg6xhv
wSsy5Omw6tqUuBcm7Ltb8gN6zeZM6hmJ1OB8Xgzmaj8IBTfzRsmU9ZWGoEYrh++5LvSG0TXO7l9x
ryDQJiD/N4y/uS7ps+vWVNasmi2FR/+XLT5/EM4fNs9ySlINcFWwaFminwzAQMy9xav2dgd6mGU6
d2RfSti8ziZLfqOWrxpkIoMetKgk6PwALx0Hl50dBjGoec51/2CaG3TKNr83pR+InMKwiGRSCpcN
3TiOaXzQHnwKj98x584YtCZ7uUnMfEu3ThCaEcJy61/BKMDU2GbXOBr814/q1BtYoEKTokVz2EIK
GlW51d8HeLZ6EqRX7waS0t1Ask0PBfJmubcjP8hTZxEY8rLiSoxreW1deSNl7KLK8zIfMVQnGxVW
Gm7yUbUT245bMU36BQIb3K4hyD0bGRNAScLLmq1AO+uxC6JCHIQRi57A2WT4R7DQ+fWvaskbmSS+
qYxcJau5212TIYoies6nQJy+2aJ+l5outknY5n7+yBEzkdaVVeYtfoYvAJQeFowqSqPkzL9iVp3E
XuHGnOQKaHAtnVinAKKNSWdGrsET+nqWMKEMZN8JmokTUOrK7/SL/OBx2VQwmRIpD03BxNW4aiK6
vK2olkJdm6BEU0C8P3XVzgseZhsXpFw+OzVsFlCeRUF/z7cPh8P3kFoQo4BzW/WZB2TGK9tahajX
VN9iy1S24lRQfyMR3FBJ5u1OlymTLyhB+Qv7UhSULq4bZH0chrzm7vOp1Unp/gqwhreW0v5nlA6J
TU7vDei+mkYX7MfYewr1Fm57Ndb0/HMVj2hrl/omUfJnX2ZYS9MYeozOkYF/DYsk+z9DHXKVZqXX
GG5qkTLAdlHZMiuCdLgkNFkf/FthIL7rTecWA7S5RlZk2aweJ/PpTFTYbCrtcSlciS/fw5bsqCmH
DVtkAhVSdtKwEsDIHfoAMHD7TzQVX2NkgIiJ1AFEkGRXN4BtFEPZ+p/Hh+/g162d25Q2SrlZRhFM
OEL4LAHYg5A0VTwgC7F6RIFft7NZNNYxTJ4R25qCodWALBg/fiv091FQdE0sQ2YATSgAEcpPLPlD
aRAcfV0wNdNQS6X3LAOfObCn7Nw0XljpBQcDIU0MM++H8gPUzD/3hohkhlCpRFe5c8IQ3B2ZFruN
WAMhvbWEWjEl202uZUQ7vU5h48+ZhqPxM4+SL4ynJSb18mT+Vlfp1AIKtvIYKWLnFN9o9xiQlX5M
GifQSkeYMKNJywIkMLPqvpJZbwObQUG+YxSO6POZYm/07s6a2eB3RPN80hfukNKQNfbh4tXo82Yp
gNVxCjCC55JBXwPVKHaf1XAU/V82Th2Z9N3MsH5iQtZ0xPj9B0zTfoVJbNTHv5Mj0Res9RJbKVI2
A4WQwCr4+SxQSI+l+wE0cJ0wLXYEWz5MqTV45+jyu9G4lb0xytUJjQhD/S5bd0DYI2uQ+w8craOS
aiLqqhQTTcEWM1KYk1RlHUdHv4HkRkJkocftWbIxXXIQw0yeXEFgCqhWjvv+R1nbwUdkTtQ4vLhL
vfAAzosTUELuAhObfLzRQ4mXYp2hB0yz7fI/y7amN38xtKwtNNxzqOuBklyteuG9031QXgM+845S
S3OHhNpaFbIkoNcOohenVzytLB3XsIpiw+I+kfe6rf5EhNBPOl6IC7gfNlT8psGyXSOQ05Ng1Q+P
yFKqsFuSyqoDnQwiIaehKGgl1fem44LzLPH6okRTwEbcwdKOh2hmJRgYJDj5ugb7y80y/3xArkGA
WBC3KyLQ6Kx/8CUsU+FLwxlcRAWRKcA2oK4ecEIRnTaQLNQd70wjIfchppeO1Ey8/o8gPG2XfK3w
AVOhG6R3xWZzIjQ9eWSKfVTHfWmgr6FBRiUnGRUn/Mez+IPgJ9B8/Lc+e6Y8iDbSOrMdb2srzrcg
oCyLDhmfK3fLjQEx40OMbv0+HwSkVk9kqhqSoaKJmTbzwtMTG+ozVhM1qm7t8cJE+O6Dv693L5HQ
BamleSJu3h/2cu+2p2h8vdcdMKu6rwq8H+7U3hI4QQ55H9H8+3q5U6I2sKdf2FTA4npNzGI6ORYh
JsRwUxHH3UUWihENgz94rm3OcaVXM0zMmREM4euermq0IulSh48ZUs8Ioxwk23BkfYxtlTvaZouO
1FdCaX2rStjOrZ+tO9RU7kYE6O5zyKUWI2qKvp4gzd9PRQ6fytsgUpKKgOUEh3FibaQ9/8mH/Dgt
Ll0PtYll7fG3MKnx5ImaIswD3idDQuoJOHjB84cb6PKw6kT/3RaxKzYI7Jz706YG1tgXF65kQPWX
OnFOzjm7a8lAVAds4i4iFlPAV5JLkRSV0yxhG0yYLxgRwrFW7dPfV08M5biJ1maXGoHwOHKShJlW
WXxrBdyG/q2/UjUHjOkQoe/2ZEI8rVm6orxcM9pbYf+61fZ1s/x3grxgPa76B245SIrsUk7ZoFLg
mlOMIgHtin1xLLLgzt8mQXfuwjKu46YdShq3+bkhrIGjxpVqknMHRig1KKNeC9UffqJLeOZwiUXv
dQA8aVWxuJRhgGXHK7yfpLbuDPQuJe02tN6Cco/n15Ap9b0cgRKFFVg0PHXN0oXd8OgLaZFwgH2L
mh6rz9CmrW4shMLLitnydFsJ8jk+YNW+Z3XKhHrpzK0RW78Le5D8denXq9HOFIPGvGuJ1kq4DO4m
m07D994fOZja2O0qLV7Fz7RLfY6K/Z91ObC187kdC/qeA+todbRYAFLbq7V4iwZzzw/4F0BFEPRN
MawxLdm87ZprcAQv+N5RyDfr6LV5uBqWqln9xHWLrXIdssr/8hLo9pbVWKAcSOZ845Z1NUw3Y/sU
u4KzPjUl9B1xEjs4+mzNwIHJqvx8EzaksDo/JRBf3LPluu1VAjm5fdOWeaZNLuknheif8LTZdPCn
TLeLNgRzUpg/LrrGbM1YqWkgvLdXcqtYI+MCC/7NqSK/gOvFFvLrppxm47f3pQ/ods1ZCjFdfqxa
BE4FvianT14IGOyz3lXcGDCWcJ27wW93aFlJrX0IUS/1zw8aF7joh5AnHKMuiIsTF62knx0PrI6/
5wYyinajFzSCPhQdTFciKZWhf6r4IMzVh1ls5Fs10rqaC59Y3f+g0pEPW5MaTAD0ZtsVgSLToMKY
rezpevJMXpIFCe5sI5PnK6U+peUcwuQydpnPBerX+1SUeeap4hAxNSqNroMwY8Z36oeskSeykvUF
RjnooJVg35cxQc6OATrEh+tGyl3QEhYvwT62LfXnb1o4D+davausKAjxGgucF/z2rZw/CdCl1pRe
g3W1PyAwrfaA4Bmd3J+RfUOo5k9ERYrUiol/iT0HeZeC7UrUWl5A9X6e1B9gUzJtH9fsRah77xAZ
fwGCo9Id1c2EL3lULYBUEu1DNN/8R1TTNqwoJs3dTnfd1876fP4HD4v9+7nJATPDWs58puBXQ0gn
+yA726KJ4BiW0W7IVzY86xR/VhrRkqZA9n/wXnjBaQDniSveHOknW+JtvE8kFFTLxr0+C3QnbcVq
Re/6yDSahwbwMN2fz94uH4/Yc4qUUHbHgfbJ2N/e7ky2dTkecGnJKfIxAY9j3twT3x/3p6iIA/Ak
uJBvaMaaPwmaY6op4+ETNkF6aEGNzsix/vf7HjEnHFyQRN+NGrficQgn7ATknGDoxomF6liY3ojx
SLvJT9Ou5zBOc4ma5BTJb3h/zwJbfOY7/q8gMyRpPKQfezDx8pAd4MPbyehy+1KodxSs0+4tot3a
uZ0R+yAym8/TM61fofh9ufFW+hZo8xBl5BQ66T6GgGRRS4T0mKfaYOVBPgTzWhPmJuo6IInfG6tW
YqNTcDzuEy/GgCS+W6E2YWRrnz2hh34Zpa9VUUEyLL+MvpBuaqmWbHnMynkdPmElCs73oTwZk4I/
P6av3J7Dwg4GspTRklc+eeMQCwchSsquTsqfR6nTTb+wdpF1S1ZKViq4k0QInMjFloIg+EJ1CDeT
4SHx5vf8aNsN62Bu3Zon86xdj4kRE9r8uShYm3J1nmM+5QSDAgf9QbnV87NeruzLnloBJMLJ8WRc
zV1wliRMf4TVzQPcr4GzmgzI/eiDyhdBRzGLE8tTQWdd8UotUmt/nVxE2jXLcBK5rWxLrV9RGo6t
xAS7nXKDyHoQRDJTFtP9vN2nmmPzyQuIIgCwPvTOOMPsFzgtMiBgymTitfMuIAU3pQZPqmzPeSf5
qs5PrwHbYWM86txeuqBHDk4qIXNhmFcPwcrcn9nBAYk7m+Wj2BZlkYkKR4W8GMNAIEWORwGYQSwu
y7DRNVD3Ci26m2dEtCfGsvS9QNkZ+Def3VA1bGgEUYLF3hYB9Mo6bLcXRH8j0/ZKWUfID/wbNKip
cMzP2meMcJz4YtMclca+JToP+AcVrgn4I9X85Uxn1YyNus2u/0ph4WOfNuaCFDgw9lAsO+MKU3eQ
AURQfct+zOeMRVHKYuyO8kjd56E8pYvaU/UA+DVzIZnhB9MnHV5jNswvD6FTaUlbLE3AofdKTcAx
KESrHunM5Rv9TAo7eHQlc96oKScgOEOIksosRD5OZtLqR7fA5Eoo7plUbHx0ltiNUhOa7Sq23Cnc
EHxARf+PlNBV7svidfpga6ObNV2G2aMu+j7F8qok+8z68RzaiRXIKYWOIjDYRTI692ZprjJCGklc
rOnizHVschoRt/3mR7mW2JOoZKksUinnDfZTr0gD68YeBm947QyWMxHHJHkY7S51a3Uq9rS+fYOb
9fgbeCEcG0bKMi2rOojq2IsxWH1DLNq/iK8KXsJxzCy/8k+Kji0g5lD1/ptopvq0pI+WEg0alCZu
uOTakOxxDWFQ0dT9IHEiXoiK1B1LRn49Ti8cGEhj9fk9oCiGWV0GEHC8efu0cET2ay0QsLR2Av72
d6IyJUCIdop0RUTogM/eTZkARxq8n9K3pzwtV+9zJ/V3dOTQx4ZKDuhO74jiW8WbRnxFzVYYiMDy
y898mbfBVCnZsfjkHGgTZ8eNQW8CjrdenYF+eBJFtGm82uoeOmA66LSdxMlYPY1tC59fvpKO2GPo
WZ0THJA+qoXh27wWZ9S8bazrebbBfp/Q5MLrkEXPwiFpICFG1fsPLRWdLSDu2Ns0ZJtJ/CeIbiCR
Ca2BBPi9tSvajhux4D50FftnoV2QAveT1l9x10cOY/Pn+moC2u/isbGLGl301zttw12t/wiDe9oT
++6WGHOHCzvQWRs8Yjq20SngIVJzWj0ESZ6MwgXUrKWNbBc5jgDgxnSF8hhmlS0UsykkM0gMnXBn
+YQ5yE9TfM90RIVU6Ao5VRvu0F2Z6ilyAuJ8Wy3TcmVh5u5ndgrIMde6Wo+vJeUMZat7Jkd/CQ2n
IQqcr2cKGBK6AHPSKF6AKMfhopS0mVH7v7wIZ9HwMbjWeGxxSs8WjIaCi7pztvZhQZ2HRpU071fY
umL6SaVIZ1OS9TnDUCkyN56zN44ju7CeWAuZDBV7isVNSvs2gK9DjXthF5Uh4ziKGb/lwF7tIIdc
xNJwJ9OqdQTOeilAmghzcoYqzbhdnC/D6aVI4ef7ex1vd8wJ9AN+9ucahTp63uMbKnrSysZvbaK6
2wPRuV9HlJDo0fTPG5xlEzFZJmRFzxojTp/fpgTtREEbAi9dxpdn91ylNA9C1TfDQvV5TRKcLBqN
rGxHLTVrcJ+03NqDTCCpiJIhFWo9UZchdcbxH13Ic4kQHIn2YuqjgchO4OwTznieiHxpv8Y79lsd
hJ+NjIueGnexGuM457C7kq6TGWpvSdshL3d5OakNesEzcjVgsa6kxd0g938Y93klJUhFdUUO0myz
AGyhqkLo+aScuPPxmVrEeFP+rpOLxrOvuhKlKoBcglWdTnG1WMnRunYw0EQj/yJJmtm7uMcp+jIq
Ruqko8dzKqQdub+LdwSeCZMT3DzcdefidMCzufDm2W/y9ezvp3mDIwjA2Rjnpaymt5CmZxqlpLUF
ndodCEUZiHwAy5tpKUEK5zWIDLWSgS3D7ONtqKr/RjLkXcybBkG7zjcF6cWnABJO3htAIf6xcq7E
CAYYstxDIU2hm2jythZ5yGRNmSVZU9tBPQAxaZyIRYtVvV/6VbKtr5J1/HZ1AEAO4PX4Q+8YLeHT
Noa3ymmqi85ioZQp5CeQ6RA+hmilbOA9aukn9tASGtDrKu1sWOxq985vq9Bx/50kCYG4IGknzaxq
bIG4pSpqL9YsuJqyHYKKAet/veTFNHSN57FTwKqHUU/kxgRqwnkANnHUvJAtW4BphCEy4YUk96TV
XU9+Nke6lj39F9nEJ7kNmf5ZiByTnUpj1Vb/K3qcjqTxmuys+djXo3YTLIGTEO2z8+6Crj/LVX8u
axyoW0VaYbSr8YMv4KFP16/ZDiuz4ZF2Zd714Ioe5RXUQHbpSTPcXfDLjrzenTQLXB297UVv4P90
RdjxKbsVmqyP9VCCVrhglu6KDoCjfB7NerC4NVoYpjxI5nEaNIc6oZfESLZjAUatzGxa+k1FG2Cj
UYL39T/UM/8FY88T315MnvKmCesbCC/XkSh2zFz7b3E1A0yNAmVi4pTPXVvzIopBUxkyxQXH6iKa
m15lzy7hM/XBZWw/Ab5S1QXg1kkExGa46G3kat6GJb9kKGN0RXpO1DGLk2k4q/xMroSvaqFt09Qy
NTcNGnm9rtYYUxMtn/UZZ5b7IYPK/ySNcgrZAzntym5YS9+db5S87mndPakZR38JdCnVmT4EO7c7
7up9uJU6coJL420iWpq7mfol3bHWIKxgbWbS7SLdH7yG2i0BdUjHKkXDqCx5R6Amkvp/Z480ZOuJ
XYsvG+NQpTPR9/IXRhro0AYpo9B5uNJaY3C5qaEyASCtJoDRN7OMpnUepmkEMbK6QsJo019mEJAF
xYCcMIQCV/EPuiob5+bUQotbWlpxfSN/Iu9Y8YNtvFCO72OKR+Fh6ogQ6uGv20imUnwKOSTi3dlV
TdQ1u4uS3ZYT5bfbAcIoxLivXI9dIjTdCMs00NTi5aSXr4ikkiBxT/XLu8j5V12iLUKpa715g88R
xQmI0YYybGAEH/l5UPpzl/UL6MHUIeXgo+yiurWICI0ye8D5lgjbp+Bs1XRMdFpA5ywP31KRPW4a
InfLIGghOg8mYsX37Jrk0ja1lNW6WqpHkUgJ0HvWEtxvnheGGJ2Gle9dD93enPqjvv6w/ovbcD3G
uIhLUGzsmk6djCuYRbaRp3rEKCfHK/0KWWLFPuJoE6s09j1UmeWa/o3wtDMka8geLQ8Vl5F2+tfK
XnYQZRGa+fL7gT6xaiq7ikG9ILg18jmnF6jEB6vgfJuyjR5g75oaM+S1w4/j6frnOxZ9BiDMkt8w
vRyviQTG5PXfCpu4spAOCfO6t+5wNLM53oLvc4+3acS1CVUvC7T2VsoHtMd6VkyZRE3Y4PqOgAvk
N5QXZ4vAmZo1s388MwCushhxfLPi8JItsS1/GJ3Qm6VGoKa4WpX6pe8t7NVO6ePeDhJDu+LUliAY
1eIPMUCwVyZhye4F64Xz29DsvSaYZTyLVfVM+D03/I7dp+eE7fOGj6nPuKWZ+5vEzIcMKY9t3y/D
SIeDzULbSbxzkRBccjML0st3IBFhR/FiQK6VyK6iiqX3/0bBWS9tOj7L4y+D+o8X/HiapGeWp3GI
rPTTx48mD9pzQdv6bJ7LLUOmTs4CG/8xppUokXg+tKhh4Vtqb1YdlM40fT42rRE06JTrMEmsl4lP
z0NHdONDGRj6y2yAZLSbAqyfPwp+5nBqGAlCE5YalSbTEfovMDEK6lXWspBHUUF+nZLf6c6+00sD
58iOPrAVxmdAIImYIzz3BXXBtss9hAECTKLK5ybq79hmrq5EC2zVFM/2qxUzvGiQUgVY1IxhrCij
+OKi+jZp7EaFBCRGDQunty4crcffBUAqwt5ulCQcX32XKTp/7oG210IIAotm1RMrGlZUE4k1ZUYT
zEjz0oYQF3rp0+ApfBeT1QPK3hE72EUVYx5djXxfGoa77SJUN6frrayOABCpKbSMUuZ8i8Sd4z+F
c4dmfbK0o721ZVuODQSLIAGuPmieJWkk1av8OwEaDLMYOli0WCo5vJhHzStEd9rGJzmx+xLxFpTa
NYC7TrUifkse/ZFlhSLzMVc6Ozvf0xzhd3Tt+zT9PlLOY9TDx8KoXFmq4HAVahVzcM37RVJrslPv
TynBUtJSdmSzON83Ql4Aib8d4XHHHK/N8jHzh/NOjP6LECyWmZfYA53dOFZ9mb9p6zFHUmZLzfuP
T1uPhgzQjT33Xkt90wgjFQ6Xhkr0oWCplNkT5ueFY8a7xhVYTAuSQ09fU3gTwt3pFFNxzLcnXjf0
3Jcl9YoNZqvjUFckGF/oVYdxhi4fKQ4jeImO290JNP6qWqAoTR/DPQTcvuXzPPIaNIt4aMUHjgLQ
sbu/QoHFKFpKOkHvyU9QNDrzIJpgU8rQHokIizZSg3n0pcYsKtGsAyaUkYtrYrLjBPQRMGyJyI0N
6EwMY3EevPcc4Dz2XpEy0YqE+4H5kw3vPSRn4Cf4FNc6WvT0rlUS0QNPJYlxEH+2IzqbAhtaiqLU
gF7O10tIT0kracg1cJhNAnHJMK5m/Kbgd8t5FhoJvXFfn7BpPj3s1cB+nUxBL9iSxnkLFz9iX5Jn
MlQur29JhDEQl5BUBjVDUTGggD2Tp5Kmld9xomBKVLWe4MtA/OQu0aPvbgGAMylqkRthy0bca82p
s+50Qj3ZVyUKX77H1k6Z/dH4UVwi2SYKI5ZUV+j6WPcl4fYaHWMbnC/nyaZRmYq+NJuS56Zopfnh
+tpYezrISGR0zDSw1nXEygrk7Lx40uE5zCp7pETY72geLIQvXAxkU+yWPXECni3iQPC8/LTKeZTB
VhRKcvFF4Wh31YXafBtjTeYd64MB3Inv3oUQfX1JUdslG0j+0RiEd8WHt32enabvOuNo7HPEZkJ4
BbrqN/QzzgQdXQKUGaEgQrZsZDC5BKHllhrN7THogG8LmkHyn+bto0bzjZWX03ndI7j0S9glCVHo
TbrgpEFeMXvwSh3+83lmBOBYc+Z/cYS5MxXqE/QxwZ+/y1iMD/Cdzflav1jwwOd4cdRbUpWUX2sC
vKqXZTRu2ucUUZL50VcGn7V67eDTCfMPJtWodasEPka4NbPFCFX08JHF6gVEk9tsuOLIFj7jRwQv
ERQAzEeYpMshEFLxk3xECAtGICq4Sa095Lr3uOF3ag+TyB/RojJm5ZJ5tVRV/StpcBzqxr6n+X8h
Obwdhz19TV0X1G7c5CHJHxbEmzM4WCrzvZOjMjDOKhlznudEzXNm0eEA74MhjkdnNijm/+9xHYaC
XgMAOvx1G+uMAVh0Mw/LRnum1eeuujvL7SUAssZsb2km4Ec3SbQW8AaWiNiNPwjPVUCyJprjdlQC
gNK8AxItYME0JGW5uHwOglK7k9Gzf4gPergK9kf6cITjVbU2gBkujZGRd6SQlmaAXVS8znX9DzY1
yACC8xaC8T/WqTwqFN3anAul1ft/fYIIYUyonnlAwRfzb7lUeZVtWHGkFR+Jb7VE2hCPeH8T2b+K
auvUTyJdT6cmgCMscz35NrTN5KkkvyJIFIw690H9DicuddWItNW3gOrIvJa+sUHV+PZFdl2NOlFN
z+HAwIkewyRzphVjXioekn4eNMPgP1chvo9tiOEtNqc455lFCmxPZNIs5j2JOd0IWh73GWgggUh9
gBnjGFdozAIgBZpXBpnV8YTVIE58B8Kte7UJiafKPhYtQm5o125MIdDGvDu3O0dRabg2iPmDFeOs
bcFd4eUYi2SK6myuGEqJk1CfODEKyzqMYfZcqcZFPspmO/OEjUYaJV1WeOKMo9QnVxq3I4lAWQsl
BNY4P7epQtMtfV/vYEV+HaTdfXlPeCeb+Ut+Wy0bLKLvSDz+Ft1nzUm1YdFU+JP1xizt7zSgTKGX
z0w1Rtduy81g0wc3YTuo6ZJDclE3wwcJZPHQ5++5QrohVHP2nlhbaAy5B3uPHua9VtyaYM3wHwXx
xsupp+QqDSNS8eseoOoxj8XadUrMCSNPgAehhdVbGsS4wuAzMzaWE8SARiUlV0M1yHLvMt2l+nUR
741GDaMP/uUu8snfVfzXcO6O7RVk6mw/LQ3mAQDv+L82zdCaJ5e7zEYyMcFrdteeea1YJ+k0Ev8n
9lXOHGkQC3uL69344I/BoFRWh/E2l44DjEWQ4H0XhQ0T6ctvufBVm/Xn8ueUjJhtzF1WdzRa8g2P
k/WxfNP5VRvd0H/+dWX+Isp8wQF0Z++fywJBBnqYZE0LyQ40EfYaSExcl3kfy9U4oznYjbDZPURG
U5IqDW3lnqHdYclxuj7YfKJaQbyRj2JCsBEr6j7faXAD63D83SGU7PnWdFcxIfXTsLrWuPVFq+VH
Cd8xdzHDr8BFtkKZwrbKiyGKbk2JUrtnLvG3790Ip11HCd53hmP2w68CPoB0XdddLOHxQkfX7A94
jXL1pkzoRUM7v6g5A9PDbgpmgE1Hs7Q7yvhWuaCyLT2h8Xw/cHE3U9qFgsRElyaRZYasBig4td3V
9jMK5337hlS0LXtC9ia5+VyWTxza7vrBGIecZCRiu5w3U55kD3axOgoA2vp6P4soly8TVjP/PyuN
l2LMyf4tD7jzZEU5Ldmpag6uEHDm0ADjxsYJ8tVlLMcAQsyrL4e6VZPFBw7zYVaMr4t34qSMMIqv
jEPCNWSFeI4NloS/jXsb1BlJrOvv97vmoidAuOOFToQCDB/n7tlzMjhU/+59DoI31OddN9t381L1
+5zhTwnf27ONLFY90rJo7KhIKSnGBG4+t6zLT84OmfG7wLpW3wLxd1oa1zJ4suSZdBoQUo2MJT67
RLxDOF4YkMMwklSvB4zyhpijZ5Kz/3Vyy19DvO6FBwvlS+OIBXTRvzxThNc0QyicXu+wWsmFJBHs
9EuHHhIjn7x5iRypRIKw5/tkfIEV2KnAVA1FdZWlMYW+vOeXSpiWfgbvUTkd/AXnpKh8AIP/jMiM
LkTGvccRJUbt360878uZ8EUpdEjjeuHm9RPW5kkaJKHYqy/buOaxANmE2uMl8acUNOmIdbULzXiw
VRk+j+1DHjfj2Wmx1kzfmzZl96jae8Xksk/8PoCsQZ+KVWLddPtY1nLzcNAwBUdRmwjt1hKzU+q0
I/xXjscPNbkJSV1ibccsTIcFwhDjjJYx2DWby6UiCn6o3BzjtJPMx0/e/uqUxc70yX85F1QCLmnf
vi5mxw3Mm+IYYpTsVYG8dY6WTBJ6F7h2m+U83utQzDBs5KfbRxmjoBBPXenCAq4biUqR0RPDGgIt
HenoSGDQ/vkinDQ6jCAX2XpW/HwEJCkmrBzeRdhzgCFq0ULBmDmUsb6fhiEI9GSF188V8ibDOYhW
9ozL4fZpmHl1QlyyajWlZYz9MkHHU0nKN+X5k0qY0MdGxQ3QI9FJDSQhTncL9wjMqkdHeQ+XUo6/
Jt7lXU8iolwL8AxIPfTux0l8ITvJXP7Bk1irwKRBwRPoAYT5NeFWytXQSH9KbKG3+Tf037DLIpaL
H10mzN8G3h9mWbkjDnJP9WKg+5vBhKnQ/GOlRVyp+QBPUrwdGQt7ajJ8ydQFl05JixXuZP4pJ9g5
XlBXYvcYRqULz+CSeEazByje50MPw3bgA6ASruTbpPdUoO+nzBblRa47cNhNaHkylM0jHjNI7X0E
HZ4OpV0T/lNCSEnC0FipzCx/1+0zvZiJzR7kRUfeK0mdD6WLYvGf8CYspyWr4eoDiqGOg5DT30fv
4jUylStCtMx9zTRBM7DMk6VFATEJFd0LpE3aViKAy3AKrD3IW0xk5HRNJzJCKbsLj96t7VrDqQr+
3RDmsNmDZrwl4jlizHdreDJFBoWpAOPd8Vq9KAMwmJFG2jOEMKYU8LXalxXf2q2WlOsKi6iyTP3F
wvTWbhq9GOPeuRiyNpkMFF0L6B8b1gaKMxIH/b2mFJgv32G4Em18JvIsZ3q3QvKtuLc1tq/0Pjs+
oeyTZydZ/u6ZHHq/Vh/RBG6qA+Zf1/qQJBQAlflLMNTTrwHiIdKNesIaeIJSnmWtXWewuZ+joYyO
uvvzxs8SvkKTJ5g7jGqCtVJnBP01f4Fvq7pvffx4iMjASUDHf6w6pTzCXS3bnVxk7X2eX1mSZery
+82t8+RV5aya40UlxPJAoRD1EWBzkD5YX+EgF8SnY6dnbOmm+S42KuoEKZ1zbhslV7jpa8/i/JOh
58UPArH8ck+Mqfz8bRA7sCxiiB1eHszCLCecQzi8+fxu0rWRU5TcAij704NSd8t01ZZKQIkUQuR4
trNu6XA17Yk6MYUcz7QsEwMcPe2uDIRfncL7ApwHpnv6bzeXyLbLZH+0/iBmlQzyu240O+PKz+Ts
/T2T6sBvcuDC4O11/UYgdSF29QoroR5gZefH8lGl/YKwsJMRey17be72JQiO3icAvoujp2kSx55h
FucvEd4UBf9CMD79gjLH/DHzNy+u4KdwaDxVtmhg71lV0nx695qIYMpuCK1izqkMbZhwWTfhEm3S
1EtRFWKFko4wmjaSSYjmcDf+XCMybYkBX+mdIUp/TJDr4sdtkjfDBdtLh0sO4l4V/7sLkrCZMQ8o
ym3HlEBrLcajNVX9+7/qcCbw/VxW1aGrZuG31HYaEHFI7+2x2Xqh8CgPaF2+fbeDwbTCI0T+g05T
+Ox8ahOZno8PCidLWTvwkPB8KkXeL8Oo4vINoMMz4P4/U8NseODk9SWMQrfc770N+OKESCSLoxZ2
C6DPbShHIftzkTjyzgX/kVO3UQO95gl1DQRmwxV326eV+viYmQ2AAp80xYmwip1PqLNvkfVL3Itc
6PC8y5/SYZiYJJ1oQmRvLdwXK9uEl/lyxHGYWHV6Rs8WaoQ6BYJImlsGPgvdPTq1kwTzaJ4lzsV9
+YFEgsA2WJsBia1uEFUoPFvy0H6N5T+Qm1MaicvYNRyYAOeawZ3p/qalGHQ000HzPY61uZhE2Xkf
wNqbjR7d4HQOyNucxRwyeEjkpnEGKNEMnkq1JU0Jq4A1rXVsKZGG/4c9WnDj/RWhhKHC1WrUqBBD
ZJ4MdTB1YwuaA2+9+ZQdA0VQN1qEF8q2ur2stPUSXUH2/AAhYKZIWaFk7YpKbmRP0x64jh47DFcu
wQp35hP89YgI0lvlZ9qch6e3EJ9aUThYobc1krBEnm6/GVkyMxIE2UISUs7LNYoKUGXMlBF8/pZu
KKE87e4t3DrGorTlrcz+lE5Cc8lcMwdQd4eUbRqkARKrsEqTTRTUElwJb5YyAmqfoE3mnzSxZ48+
LreZ5hNrbw/JqdNpqZ2HRkv+FIS/vFgArYaxfqjfzIS2uFil8jrH0hf0a82fkq2cTKCTajZQPNeK
667GV3S9j0cYD+xAeFWVDpCA21sp9gjUHF88LbePhTkyDd8q65xeVB7iU3WQjRT0VYXsND+VHifJ
gfXweUOiWy+dKKkyIiwgprnQNUmpjSWR8fc9IvF/K5KtfwWzp8Pj1xARGZsQNiOPbjiDaoK0zrSx
dVKi1PvVBqRf/on5/XRiiYE6gjzZnfH2dhwYj9xNg/JI4WA7USxgPcQvZHznTKQWpdtONU/CSjjw
VJr2WUkc0CQVT4H5Y1m3zuChWSC2WZ3vqZ0s+S5duMZ+9j6qlIuDiRwpSgwuAu6lu50jT7YUZRov
7wybXOzvN5sSKeSsGcvIW1HT3hFriiBKoKCTI8ijYAHykRnJALwMzI+lUELz0f9jVzK/h2ELk7gU
hUxFLOqL4fj3leXpI+fQ21MVlNnFu3nAKfH0hCKAJf44ujWVZfzUr/74Duz9TFuhcWJNtnIGphnK
Lqap2bkUvBQVqEAbG3szUbc24XJiEK/c48sqr4zts0/8yr80e0LrMo/FWwB8g9DfhYHFCvognflC
F6qTXki/QDAOaKMCYsMcQPf/vJJIGdHL+8hMzT1Lcdik2RdiiQQa5lTNzwyStlWcpMDXcUCPo3/m
RGdkTgUjICgeDYx3FU+SBlbXVBGGQj/w2nqLHW2ZDefPycNS3gmy5CxStufIwbZGZP2JuCI1owA7
hH2hO+xxtZoZ8LlTAk/nRGfNNaJcNDJhX7G7SddF5WsZPUglyNLNp9hACnaxOkRCw4nJ7dPdecHQ
LQD/+rNFoQpsLV6jr9bDkyu8OY8mwgCQPdRoc9iagKNFym9fal7/rf2R1cvcsfFvmiLgSadNBD5p
GVHnaUaygvf7VNgGMURwJ+8SbwFvYnpx57FcXnKlHvo5PrXQLV5dZrrqmDVCGQSv/Qa2Lq/T/+dX
+hr/22LWy9dsLqi/zyyP51PU1FJtGGr44R7NYAmYdffi2t4v2UJLTvKO/7l7CVfDKtuNnLOmk/7j
2dWfjlIiPYVXSORL/+GEkH2h7drfATMc6G5CoU6++7DXPQzWajnJv0sx9+CuUT0PyHHDy+VAxKhV
N72v4a6bp5aX74i6huF4+ZhXtRu7NQ/iVU9zLhzF7V2FBkI+NGSfYf7rPqF3NMaSxZnvaAMWtwNP
g7I5cDzXCr16J/o/wlRivcoGyTVp2kdwbI5J/UyXDEMH+W+15+SVDbuw7b+nWDK71XomsGUp5YUC
fwzi4NXWu5F2LlUPRvLJJ/roaY3SkLf87rM/VpNpGRknpvsikYXKrSlZ0F/PRf1zrPrusmavpKMi
Zq7l8EqYkfWy8XSqtSLT2uWrfyBhAusui9OwREYmHwFXEw4FGJ01Oa4hsrU5lDwCKdcKH0CqOoeN
NERnDH5AMB/33LYg+yZ77BbFsXxhm16mOvrn3rVC+u/4tmq5Kw6RhIPoj9CEPd7Dr7sQ1dScOiVU
j+lr7QP25wuBaAqVa44tkeRp/BxUdIGdbXavj2bhYN8SR6FkZbuAsVbWtfaGoV+HR8TQ15ncqXRX
1xoujAUaV/KrlNhKJRwroq8E+TrUHmmWN+r3tlkHFGAG2OwthlqWGJMrZAJgL/PGBAhKh9ep2hQ2
tpoP2rHa8o7Nts62Od51shiHRIvWGN13BICEM6xElrN1xpGLpizuWvPRAyFQZBYi25/5m3vZOeUB
sU+70lMmmTQSp/nuOLcMdzFnhWaHZhKQdLyTB3pYjTmi4yOcclNEeuAjdPrHgK8X5mC0TdLDHB8V
ERYMtv4jgoSKY5CAsnCJTiL2pWofnmWQa33m32BFEG1pRL7Ujn/xK9t0iJ/5NH/cs59qYzFWlfqO
wqfL5KR908noSdvPCWBOiQ8qqYwZSAWcE2SI02MrZKsjkwNwWfKb9Lao36W97/qPZd1kuZsI57sx
74TSskqWYDZSxVElbZXoCVvYUVk6J9Rlxp5kpU8ElzjaUjdpCoCShG7HT5ly90rJX0Hf6JQUaaFh
S5jNCgpfSjG2lBMPZtqVliW5+OMYcr1rTsMGr5gDukmxDDQMJBVo26BrAAF7/ByThW06IVwG/0Dr
QiXK3BWLF9CLtc7NG1gPBu8qOI+9isj8CW7d26EG1uGGzHQ3PJGAAhpfCGR/nWfNVR2iObYzbixq
Rw+nZKCCpXaiRMMZy2lOZFIqbUgTcply0VygRK9DlrF8S4uBO/B9lK8tkqA+wtYXAtedSoFeMpGt
d4Xx/M1h9Ei15cktA2bzNAP5D/2r1OUeuMcA1Uv/Kv2CzJeUSKmjBSsz0+fQIWBijldmaIbCX/w4
EKRyLVrQbGdlIE2qga9Iz8w4qPUeIVC1kYBOGeLF/nfTG5EY3xtGso29sQmUKZzDRIIcXZ1JILpb
QhQlv8qHoPfY+l5ijtzzuSVO3sHIchVSzXJx1+o7AbnL438fyE71WsYUtapVc63OPXuBv7Am96O2
t2R1NT1sYDHf91OUV03mhopmWQjIBSfXMusvVsGvxl9/Y1F+6EGmW7L4Pbb5SnFCAbVAOF7uciss
JlCGgtVGrwrJnRUz63zw0jOZ3RIuRSz8HmZekRc9bf/1sulHeiBPgJcSofsHf64bk3OPFZeF0G9p
4jkWgCxyt3ysmu4XpseSWOPLdwP5f2gcm0SdpHOIoKgYpEP0v+GOp/7360tbSuSTYgr1YaFy9N92
R7Mt7BFJN9um1tSZVC8Rbv/l4bmm0KIadOWeAaFIjtInD0TSnIqRVdVP1LQM2yp6FEM+gg5rFAeL
Wexrj1I5XGZxB1Z1I0I9LGpvo/Zp7ZODdTu3grObTBwhKZF/mYkvrWbGwZwsGMo+8e0Ip+lymBui
DIi4FSnQ2BJflmcA2iKcrWNb/MhhAMBlTSIeg2GYgFjsBAqXKI4LsEjfVA3MOuX8SAVt1N6fqdAS
5g1MzbcplbmBRERMzFDVzPgn76v5BLtZsI+AYGLxcX+UxFeeGaYjQAejV4/9o345VOR70sX+2Evp
hqvEPuGoy6irysdlVf0vjhx32blGeLCzXCSDr9fj3+H+1zGUhW9vjQiSiYMCgwHQRI/ZWds6Q3YU
phO0WA0BLWP8GPkQlr8rjOs49PSY/RuzcPAFzrGh60mv0bze35SMtqesSQxLKcbi1yZvqF9XZbHD
JSR6T9UPNHJPG0w8uGJg8NjUzjJuln4hVuOsdMTv01qavcmGjSY+rbyVe39/MZy6DChl6qNiR2fr
8TeWAoclZamok0UaQJBTxBvbrZWOM/utwq9A+OMFO98LQdCJGaus8nGMcW3Fy7QESlLOrL8V59Jb
lc+16STaEcQ2xGGUD99oWZsIdEaKk9fYQ7G84fKSea7bAxIw9CNkl842qzX0VjmBFD08z1J2vHWK
jjWy05af++KdtSD1XB+VJmXVZLBwSRDh6Wz5X66n/kW7d9WEfkqUUxFare77gNzD0aumV38cuGD6
vYNFTlXaCLzni4v2IDrH1EbuqPhayUKOuJbKGr8eInRpKraE73gMVg6N6W3Y0z5kGWIJXyFiixEW
UO+yir+anKUytl3Nb8OcpONZjH291i0A/yeCWY2yCQKUQuhsFnUaBPHHlCDrGhKSEQyklnr/76dH
HHme3/4iuTaWExySRB/UkHbBNYwLyeZLgX9CltJ3iUeGxsbEfePHydtBF2XsVu9A/4yhPeSrmeQb
HE+HZdycJKaE2+xqgN2/PbQEuxeuoj6xj5q0MZlLhzlOLuu0JWb5umruP4pTq4cUEjIMhGvHLceC
Vg55qT327PvuBY0nPX4RLg3eG26KTk6QiSW7aMHnI7zgJ6pVpp2LAVescoita8sgOGiN4EJAxIvd
oVQSJbEUDXSCr7pk/8StVMg14h+48eBInOaQ66ByluH8QiSUmpUoTbz15dZnfn+A3uYPrem9d/Yn
unNtK3FbmmOfapuPn2JuqMxIx0fhLdqKPAYwj8cpNrz2oEB6+QcJrpnAEqwXnj4nM4OTD8UTpqon
knlmPAyRmUknYnj3S+9GEwmtChDmQAvEsm/g1l4y0lBTdUq+0xttRfstf9Wo2rmJ1gzw/AoE0I8K
P2b8fyz5pYPsiqLoMF4U3N0obrgkcssOiPp11L62KODvcZOdO+C6GMXNZGRJD8vxxc13m3NiU6qO
idZztDJh+MRvFhMQrimDlL8nuwsCAlQKYFSUzHraQYKiJlYWgVd+LIkbWYQ6qoCDk1MXSBbKPeEW
vHQdG24I1IvZsussvyzfvV4nX/UU9wsuBWQ1eU1PerTJNgTy6BsHjuddwuKBbcUelMStEos5FLrX
J/JF/mMU5h/CpJlg/RjRlWAs8QompbHCeV7JFO8anBead3eYIg4yIRHLlPruLO2NAXXMysMph9ik
+ApU/CbD+ut5RJGMPqGdOGBFX6LVitMBfg6Dvfq35kXXIbkw9Smyc4eHolYAD+VclWM9+RvcY9o8
1wEX6pL547BZu3KKNKW28MJ1bn52hAlcVp7JOnvcCIwLY/PZqapHF839Tlf1zWwzNOXZgcSSijwX
HwkufEneDFM8XuXJte1OlXygdwmGz+hKtEk7IrR98aWn0HL/YBp86N5hqO0VcyhIwnxTR16e6Jkb
BgEEIojmq+kO+d13eD9HKIhMwbdPS1MwxCBhjk4gCvJL4SGD61Ab25k/bs+XxVOveEiYRq6wcAnX
pP1EFN6fZyuIehQqimudS31bfXYHC5JFNpOZln6llS+ausIzGminDZ7GIoEkN07W0PR4CS+oyjP/
/DyCjHZcOuP1H/ho/dqqtDSENVULTwIG0ixmh5ZBWX8N9L4n7V0JWZzWpIiHQsQgnoKmcdKiA0qF
bScewkKUPfLyBEDF2RRrHNSe8PUywU8S2vo89+ckC9DTqbNlHZuzSxGr9yU25a4XQfGczuFtcRrK
/rSk5YAR37+P9Dv9bQjU6yKndjraWbp4Kux1QHEj4zQjxTetAFy+j+JYcwSpV2LtxmKvJDzYhjW6
/1Dz59NDSagQv6Cyc9jXTdGvu6DfxfSN/tZLzZzVOpQXqNpRJL8M6f/EEP6k1fQ+Y2MVmN5F4fRk
EiRssQK9Ic9NeHWj7DcWS+MPeWcq+uOpuM/aVPYCW/uD/GzL853K+Nf+K0krWThYPDLzbQC3FEQR
jBi8eW169yAiyESCbWnXwWHJDmDOyHoNqtKKCgvtx5DSLo31JtqBNzWDTcC43g9RbD3Sp0QeE6Nu
06AkoSrvvwmxdvulntksbRGs/eVKQmGGwsMTYKzLwfuiuRN7yR6JEv3FYfaHYgL4IHs7ERyt3no6
Gtl3fyIgz6CfW3l4mZjZMl/OJgvn5AhR7Rfk15WLdNGkJornZgedHEdTN7srXWAd5Pq3LkgSSvnp
l7VJmA4aejvf51sJgSrpXSvy40JQniOR226obYu6aaLRq0a4Qxzr8jGCisMbAN6x6nNByX9jbaIq
x75ALGSQbWmC0e/qAj8XY2TPdFF5fTtJKKhByrpg/6i9jzUxmXjObTHeq1gsTLwKlKZs8YekLqrv
e80zel7koXz0c7WxYvCooTaCmX018zC+BL5l3EgvZEtWKTTvDA0qISZg1FfuM46YYlcVCFKM+Ql5
gMK1BsjWHB48dH7W0bbultJtaXuu/zaWZNN5IhUdomW368yZRg6vKQ5y9SdY+rNdll0w9J9YlF4/
XhQG94Req26L2IiQuW9+yQG/xixYh20wDW73tw6BJ0xBsbccda/D+8qrl6CeHgswuPJhSVGXMy8C
xIZsfk3QPIB4T8TkV92IX0PNXE87aaKV5+9U2axToulst2X9fjcQe3ZCT3hb/0HvoOw7Yz42mPk5
968s2hqoksjJb/VkRPPHjQIgdRRAEu8kGiMD6nqjSxVYGthOwa/0Uzao3lR8abl6zMqnmS4JqESp
4g4POsvN2jRo7jJ/na7H3sN8vh0ZvZfBZiSsJ0/2DqOMqcvPxXkLZelE7wXzZG3pdfx6sPZocFEO
XDlEFnZpc/FDSt9JdFXVlKKe1Le8OoyhJh9TiHJnUz1H6OlUzsvAO35BGHmcBeiVA7FGlcWOIlXH
rvQE8vydJGC3cXIhC8LYRH+AoqN+8TdCVJG4a4SjhTGqZvBEEhx7NPtJxOlf3T1XXwX+GQ9F4jHe
/JbJeMK+fWoX+mTgrCz3uDWJyVZxGUCcZgKr4pucaZ9IYvsiOmyusPufwZbojYTA29IYysqpwafz
d35nuEvyptUa/YIrZR4JmrUtXL9YdlZJtyMTkv14U+wDZxT6DtKf3c53qHoVBdE6A1HB0bnxky/K
vaeWf2ecC0VZmn4wIGmi6S/do7IWcg3/Swhtc1SPns21doTnfFMtZHNDpxrlFQXtSt5hgK8uxrMw
fGEdQGovdjvuxyofcqHCVZ3jfuQICdLTaw5oo5r9JS0lPB07OZavkZSSILS8LQBMkDlpVd8P2o53
X5fJ8rrLceC02H873pyVkzOCSV/6nbK0TlLKs44fhTRN7NBaGRIWLFlXgwPoA2BdLVY2BRTyyPAO
b/oc+BE6wEqPkjNCzQ95eUeKeFZ8Of88PQor1Ef4vORGAaiABrtOVtyTPspCklwbX2evpYORn80V
CC/9Q17GrGumC0UrM8qMirxNW+spBVUZKbAq9lnrN+g5GK7V1A5+c96BtSYm1+/f2tsE5KT1D7O/
sc2hXE8KO0WgqDyzlZMWemIdcP5IGsS/7jmBXYVfu3lezzuzRAg6tMwZ/jaXwv8Kuhi77FjZhyfD
I18lmIqoejwahjSwLrXx+BXyA1IjtRFjONWYE5Vrlqqy4riTjXRFhI9U+7cjFBdv7Fx1kbDRHj1q
Z02iuoQMWzgZicz7F3mzcy7s9rdHxte0jt2w+Mn7iUzEs/AVNiYqb+JtKXBaViVPHHH4GdlUHQTx
UeOYHYQjpqm25DhAMjwGTLruTJn/CWz8sEsvUlJ3LESPviZC5HOxQL55sF0+xiQdT8E+I9jhgmYg
oY5DqVckBaHwippF6zK2vdWWkoLuLXVBUtG0wxbeA93NgFslewdfl52zouLnVD3rx/4bk8DkeWca
G5q57IZg8rgIzF+11w1YXYHTIv+oMu/Mv++CN6JPY2vmOCGCRMcRRK0aDH1VsrDk/3xPPRLJkcMb
xvYFibGpu3ABAKa5NBxZIyXvtzZ6U748tzh+Got5sVO62keDw5It04ainJ/INMYsNS5WSPlpbsp/
XX1GqSzEqKn4CF0Op+8Z72WaJjHohvzlfKT8mqONJ4ar/ibKkfb1ZTQJbS/LYd/I63AhHxBXxHa7
evmkWea5hsJzdr8v4TO8S+ltBrssnG2FYHsYRD1M89Ya++NMMqo06Irdfk9Ye1RzIyx+ZRoYZodg
YyG/dZS/ed3JGEF76Uc3f0xKZM5qvecV4avMa/H/m51CYxTwJPwTIzke9HVB9lcLPq7MbnkuKLk0
oHZWqadOhlIoLFHgNGrMmCcnEDzKPG3shf21NOG6M73RAC0gk0fEyyuSHb+z39Tau2int5uRhwPd
nOz9Gmpqd3F9XCoLa7TozgLELb8kKOWZGnBVN4Nogcr9oNGLyDXq7ltncqKd4NbQs0FyRjEOtVdp
yYXP2VvI/eO3x9vkQDYeLBlBp7C4q/oQWkZ8prQqb5FT6GhwCPm/lM45FJK0j4YmcgE3FUsh3FuN
2g11jBBhPNuCT+/kGdzrVqKomeEH3X6R+NaI3dEMGC73bkYExC7H4IDu2aEwjLtFmSuXAHCye/0u
XOzdIrsFAYUF0mDj0mqMt6VD3RZwJ5cCVnJUNR0/3/x/6wTjaV48OUdGybmFT4ITiFv4NVc1EOgs
49Jnb24gMBLdmxRMRvzIfcxzG8TomRBM3p6W81FR/UjrOqK5ABHx4XP9LeO+hJfpJoeH4t2lpKzt
QK423TWaxrgjtZQ8TC4D/2OI7KM73SL6pYLHObQBl3maJR23zEYLvfHUjtzwY3dLT67Dac6+9nDC
YxC4JST3hNN943zlYLm5vY42zt2MaSwvEvKCH5Ml+Nz0D8uSABv4V/AwDp+8kBfakHApkEl2lGvA
n7+0phhyq95WWXuFuxl/PUTcTGqIpTB3YsN8qSJfZ+VaVpRhngAREgSTVy05KeQ/Z1W+3ab705kT
Yl7uexUOJJwQT90iRQY/IWP4M21EK0Q8e78WzOgwehKNkbJeBSEdHncTbkvMdz9uIgXYJC9Bt4uR
wSomw9n9kWf3OKwFYho5lm2P1+lPNTWeEeZAUBzth7WYQKWF+6z38hVfFraHiJLyWETBefEs5pMO
1uRXvUMff5NacxB3USsLR6owU/eNRPurj69vFYy1gB0Ah5PUAiuGM8lEiQcx8m+HW6EOEBploRmP
wtjFnk+A5kiFIgujWTk3PXoqaR6zyVHWnXEYJi64tQlR8wNl4MQNcmNu3OWzIUyKvG5u498gJe/O
VjXnM4o4pw9BhLabI10Q64ueUDzU4QzX4n9CI/R7ln1nnYNQFn7TbJQ6SJurkkj5BRMv7Ut8PGUR
wRleseLGPIbS6j1nt4zOQZmaDml0dgRhDGpt2BY1XQpFN1yo3qAwkdxZC78qSNfm+QkvbSqbRMrt
EZCpl31WSI2STeVOhYm8qaneoAO7T6PtW0oGt05HSYxHehkqmO4NP2OShU8klmH0C/xno+XH6W4I
inDY8Trao8b9XmtxmsQbwaLunRf8Dct6w+wc49H6CvzEOQufUfwhihK4rT/7GrzwrZ8M34RU2qCB
8jl6Tasd4O7LrIm+AziJkYYUZ1B+Uut1vdagcNQqMr8ttevi5+AhvXVU2MSlTvX9yEgaJHFD3/ah
tjbioy/qmOxu9Zw82EMoexzDFmJHSvJXXIqtrw9sN5p59eI65uWPk+ckrDyhEzYUzwfe1xEzs2oE
hXo1/z/gbdNCxeYXbxZV32MUp6cA6DOdKnT3mOfVlFYzRctoFLOeIbAzb/6tjO0bZsWDNl94iVkF
tRj+WxwY7JK+/JeWE9FZMz9Razsfjzt+qA2kcHXplki5ilqtzWTymetLGznT5DXyKp4jBg8WnXys
UUaiQabUwInK9MYj1D2hCyshnOtpJQ/92WRA1RV348ef/0R+zzx/fRLj5j99gIhOAWHufxqHS1GS
BIsBq7xqJH4x8HaYtDXIaP89Uzrrlb74EisQeCba3OFfdntQ0wt2X8LI5nNt1zmyUg1gWyEm/3Y/
XxDnFa4rLP4tbZwTDmk2beIZtAypdc6meavCJ94Y+OClK1AmsZFKjwyFw/L5REJSGowLE5o52TSH
7DI+XY0EENetJcWCMybTCD94HiVkQ6GYN9maPdw9Up9MVxfSEHVq4K6uZgEHeYyKr7um4IpO/Vpf
aAR6WdC5Y/JeCDoX3lCyUNc1ciX5GZe3h4vQhuu+LOFSebUBJBC3Wk8reZeM3LemIANlOb6gS+o4
4EulQ6YL80WsuF4bFvmjbO6S/906pe5c9vFyyhrLZpQyjFZUK/BU0R+HP1KhTt8f6IkNdNMkY3rV
ih2wluNKM2z05pSBRfkRKn30UmzwJVaiJZmQwOWlQxUlHDQPIPoy8FlfAf45uRo+DwvX6Ho+iSQ9
HKq2dpVzkIPTn9DQbBCRyOo6O9WsJcdke7qOcNEA613+gJlvEFn5UwtZoTLhIRxUm7tZgMFuCtCF
UpWSMINRCb/0L3vvFi3J1LIYSJr1WDHqtiV47DtdLCqRYkvveEr4TyPzrmuaEnS6P6L6G5JGtVvs
q9W657GQMlNiNemttirWVFMhO1GUIXahvHDcuHU1IsODZ7systQug40xADLqUT0vC0ajqRwDFfCQ
AI4r4RF0l9Un86unW1F9GzdOJWMtzDshiLEuIYoVt8ouBAAkjs0mDmBlv5yz+W1plnybhZ4BWr1W
5YzOPepk+asFjBkzVMZYcT1e1TaxlHmq+1fA2RvB0fj0KVwktBlIXR18+IpXP+Zb2ViULyVY46FW
VeXtv2Fo+nkSiyMn7kBybBrUaA9BIZh1/GQMQRKFpgbGE6U/L05zJAw7mqXCPBegmVGYpTW9XJ+V
1VnJELvSJxOAqhPSo7QK+PrMAEX1Te9J9A11lMTGQWzBhO1Ma8E+mfjwv8gVs8keQPZk4MP1oOeb
rD8jpTED2vaXM+lh5nUOPCmZlbwJ2OH1VEg0MH7Fidn+ud7k2UDMOfm2UnWIulLSJhkiM3Y/zNkG
sH1Vi1NCAlx6wzoIgfaW34SmGP1u4/Z6MaD1CELMlU1ai8Ik0iEF0e4Gz7jzirqb4LLlLWtzxoMd
J5fzeQcCOCymTTB9yVitsz9eOwu5rQ99zQ0a87CQ/bZ5PI/uwyQPxV/M+vSQTGiJfU6ffPR1wPa3
FADfPXknNE5L1PoJkFge1GCyZ5gLAY3Tf/fvmbJhqGxAQWT1StvWrJNVnxdVA3DsAWbZm57XcCqF
FaB+R2g/HYUN/aQXOG7Zh6qd0dFx15mwXrWGgakdWvjOZJGf+xb6g52b+30ydIgsH5rMuMFLyyr+
2VT6SaNy10YBDcLx2BB4QV2LuPnIsgBRAyiE2HdcOp1iAuPOnO9RTBBwEhpmmw9GP1xw4ibtuF/b
kkf0W02jH+Qu0/oEro2rgOo+W/KEBrDQXg9Z+akr7QoPg4M4NowKbcplr/b5KQY5PlOmIr+c7igl
r/B1w6q/5htx5/oMKUWrkGrtwlXz9uCaTQfMXuGbLDCaDI/LbJ/MPv0RxSzAiENIoae3xOjgv8Wp
vugwdLo5QIzxaAslZcEDBggLtKvcdgeaTUMzGjMm8Hg27vyTTVbwO1sEN0Fa0U/wj84jaQym5WPG
K4wv3f54QjKysbpMBJPzPqQrAu4m3J8/S1zx2qz4U/7VUUgPw7ypH0WpCjRAQ//tk6blRJfGq2Fj
NPgnjiOEaLUVbsxkss4LN73iI4stRnMEX8wvZxFUuuDMI1kXq8S3WQ8La9lOeYbDVZNYoNXwCpYC
+aQkIHiWkj0atvKHGggwYtbO2Jtsfq6DER2Nx92YAnuSUDldAzP2yhSmlf7/D4HJyn0V2lh61Qov
yMx9cAQGtyHmL1jArzAon5O96MRnFsJu3Tga1JkBJ/nuFRBHDStnt1jyJ/9eOeoky0kq0FZ2JGAD
ACNP5yfhkLOVnfj92bTQmPditW4Nc3dtVlk/VzZleZ7nJyxRqKXgeXNRPlIJgY8sGM4qMtR7Y1gC
8VUs7WWa60miBNmCEA/gz2YB4tBdeWZtw1VSWTY/Y7HE/TcoOScC9CUPsvSXzccJ263r28z55p8e
ig5Gf6iPFd8X4ZPD2nksVhl/azuIULcXA4fAZrv56KbH763WNucr2GnCWZebDHQcOABrE9S2lvD0
WL2dtq9NBjBXLvJ+nxaqAYMJEnpgOJahmPOFyXs/BCD6uw2CmEp/uFn14TsSRhjWK1bdIaG6kB1a
sT0tuTuqZiFCKATIjVAb8x60szOITk9CSJT6Oc2HstzW3zFhWRExVmRzIME5rT+PSBI23V/o5tFg
SHizkUiTZKiRT3IfXDxcCKs6V8jEhuRtnE7rSW6eXk/tumelP0UGuOpRwJMpeXtgGzYrKPioIq5Z
87ZTnOcDrqdCtYjuVrZ+hdXHeIkUPM9CF7F7vyhQbzy98TGw15LmYWPAvAtp4iD/aXpluROK+IEo
ITvOInHo37lOHRruxD96E/baWyijcISp7tj548f6ZOIUz4WpXf0ASvQEcfVGEKwVQ+0mog51Tg3a
oIjblAbkbVvFtndX3OlfK9Isrb8ElOFXgbqLqrmvO378hC/AQbF3RYmtgG/SPvKWIauilCEfWp72
IFVl+Tszz9GzbrxFAtz13rhcQFatXWY1CHfvCYu6zXJ2YlWrqeJsdMkYeHO5VcfZyJ+P35dPQTGA
AKiejmHtVPK4q1UtiiNtSWODc4HjpwDAhCt9gOzEmuVfquPID6+pYzK/0XOX0eLZx6EKxCQ70cZP
obwfmW6F62jF0p1lcsmv/lqzjR02js5guZYaJEiXRDmPCKE9cO+Dm3Avqkw7OHVxrQFUGDhQmVDM
PvvxhaIrIcilWxGrWiKA9WfrruD7hgWOns9YXOMxVBwFkJ0Xyp/exMBDtR7GZTYOCRXoafVMxYpF
QdOYeVGGTdK2Po8TXrNN4BQ1SVvDUYa0Qpgacv1pWmuttxMpJFJIoSDLYgmPNjcFOuHe62SVU+ym
LjIMU4oti8zRlmci1VHvNyoKVyk1ry1waRllwtrGYHMN26c9P8AivwmdzDuEwOmmMkWKFM2qRYwY
Py/CPSX6fREoECVyfDDYCwOG2ONg+mZYGXfgECXvdF/QnpU7GRFI/SNXMfpNiqG2TI1sJnu11KxC
+ij7YAtirE/uOVxe8JtOE18qB4Kwrwua+VwDSTMSsVTpD2THKcuPKvzdNunHmSSDI5bruVGbzmB4
rAMFb37WHPBzjWpbJc0dAb834z4ymA/UYp+cBdKnBMSxVFltp+nSiNQd6IWB/stmg6MsAt6B9T57
5JzJf6l9sf5DhyTaZYXzr3QJvyHwuPvsEZyPUjWw4dBZkeoC7btvxzggixxD3sDaYphmjjwL0f/Y
IvDKJI93Iv8bHEINI8VwdEdPVJy5lubigBinMXpYSaUwbghxChIP9UqG/Fyb1aZF4VdPePozr6II
XcAbpuyrxHBSrFpjZh0fLYNOi/lntKIymxYDFRFUeOo8OgZ3dUKEBWabJFHwBvg3xz//j2LGq+a8
wgAGNWAEySuGjp74Kvavd6f7IpVMYPvaMkk/v19nuti2BFjzvuillnQpYIEl3aXcGwL2/oCJflse
krzAb0PTGvX36Qx/fun1WEFvVlenzDPRjqFAjRG0ivBgwFI87vT3MSnQX5dJ3HhdTAZiyi/9dBz+
fTS213r/XqakmcTdbuafEbOu2LhNLHAe+ANBLf4x6/vMESQHjqACk/7qDEoCgdbjwVesLUdSZaj5
Q7zLK0c/RrNKvH2LLApOzx6B0g1lSVgu9nIcKhwNN6pN0z/asON8k8V9yE9wIZZSZ6XwfGWJ+nS7
autN1PpqUaAnrbdR4NNxBeEu8H3RVSVdUGKEC4nTIbKHSZdD4aCi6pmj7jWPGGa1Z2NBs6usFDP4
lcCcW818499aYXAZJ0GY5hdF2xkuhqH6Ccf+pXQRs2CBHRjjcq7Tn72+Qfdm3s2Pnugne+X7Mhnb
3mekwyu25rtL/C2JzY46d/DdZBQaQzlB5hmg9RoLcbrxgTS6NX85WJLT2PFVACuxpsr6CsDlSbhg
etJOVvbliUAbRvioCLfXeAYrPPwZrBo5r8s9O2le8NxTx0lbryIHei+18pHPxzMfwKSDhiwxuFQI
ofF1Jnp+7VtcQF5m2alTQY3SffBJWf+7md076inGe/3RtOOYwMNsfJ9Fz9VUzy64TljOLTJqL9YW
yRTIU+NBa4u12OkzE+ngS/zX/kWXu5iNfibtieM8yIauvqvGnVc2BX0qF7TA1/AMn1lZf1WJRBY6
Rn6Kk3CYWMBAbhL/rRpNnwtmDl0egAoNHwtp/YjdIdJXSOFOGK2W2XAq2i9SPxGWXrTlOdu3n6+/
90nvzgCes/zGWDAPhgjPHFBicuDKFDIT3wKcH38V0keJLylLX20uxJHcmba+M9gRFWfy8Af0Udm/
e4qR28F4POzcE94DxP3mlm/gXcsiou3SzkUU3NRzWBcLn5DBPOS6ggGP8Sjtfnhwc0Nn7ShACBFV
Y0Gwdz1k37pnvAGSrjMYa3s84ouwlGSDCkTMgNFti2l1lAUF+f77q1ry3u8GHLojjoKFFAmm1xp/
qCBD2tf8UePdMUXNX+eqi5cath0JNubhn2aVL3eLk54eAvpCBYezOTyl9NxXKdY8vTkTzF70gMO0
Q9kernKIkVQkKypZaPx0vdI8w0NfdKXO3z8avU9U2pEn/iS7RZgjzVK2nSG1BYVlJlWQr+MpOq2G
olnQpVuXtcfctsnt3Wz1a9JHiGZ8BoYjYVBx2T30MilDYsTUEopLLFauM3MdPuzD5Lfd0EA4iUoo
X8RITUOsvHQC+5j181o2932Q9tneVLpOluqEJeCgixeEPUmcL80jJcPNFtUixWnSaAUdn8lhNcpx
waAWCQx45mDl67v1BVTe0U4fdcvnNN8s5EnL1PN40Ofk7rO+IS/GZr3KUzLyVQl9qcrMuD6sz+PH
U6Pkqz32zI7N7QN85WTXsmX4DM1CMLjZOWo7IKTwUTO9dcDpk5tVzn6eJR3iWkocf4ekNPrmEPDT
LScIseh4zBUT9IpJ35SFvnKRb06FHcjNjoPsgVuALVL0jnBq3mxgTcJME2sYpgI+Q3Flp/2+FwDL
IyZcHbwohJWz2zzxb1cFA/Gs0g8JreJLZKqbPyh8rl/g6NQCTerTve7/bnndSY7G0Dfso1A9p2X9
E5jWiU1kpQpTJ1pT7C1/HIY2HK+UKeLI/EydJhZ38OTrjGGDv9c17o+SDrweibis36pufGSHYMzm
qPiUZjdNhakvRDOJejFJ5IX5C1Arua/NM1wXpEq8fsI/YPuvurgU0aOHZcCChZYA99bYnAdMChe6
5aFPL4Wt0YRH0DlDaJ3GAl3b+6pviUd23S8uz1hAqJLFoiwlKdT4NgrgyPl9cWagEHoGbXvfQBbj
NvsmGRCXGuZG7Q0hZI7gp/mtF2aVBeCJLitVXRDzTEx+yRr3DPqqmRpK7SDO6ICFthcaKsqQqdpZ
XZHc66kkdZ5VirT3NSBq3zo1jwjS7dxibhQTTotv55aXcVN6zBZkw+clHnmvoAhIVR1O3CZT4fsp
8TfQW7qy6vh6UaB0Lr3XUeFRNk+ls9aWtr1hS+Op+Jg6mkKwWbTMYWlaoDb3dlhgL78BRIbSNLN4
y4v27LP6CXyUwc/bAMBLrYVR/NoSBrMlFn+k2qgO11x/6px0Qjpt4SQHYLBePVJSzsDW2b0x7W32
0FUlsAOiXLEUUg3F34Kdd5tVS2oGYM1wzoJ0H3ye9V5lQjSGmFn2YaoBRU8+2eQMM2fv+q+PxGOl
9OH5LMOXGhX7l7Wxl7tuFUFYIssRJ3+O9QwkLEnLE+eCRyRtqJ6c8SMJD1IEM/0k3ZmaxAzPxHBU
Bu3vlDRVwf22wWD/SxP9SJByfL6fsg8VfZTWB8T4Yfhj7gL9AUN+pJVSjnTQ9zZ8Brb79RJBXhSz
BDeKaDXGWcOgdSLzt2lNO7RiKUpvJgrXzQ55PNRuIrS0ZLc3mRlDh/ygfGrm69meGZWkyNXz80AM
MfqEbYglNcG9PjMMsfMkPQsqOE3b1E7uQ3i4ADgAjNvk9nHsaRcDhIa4dH3GdssALfysh0UOvZnT
eaWNkpJNNlbOuQ18+I7m7fAPAI9DQYeLQW7Uy9Zc3EWMwT9r6Fb2i22tBmuJterZVr3vzlzJC3eA
0OV+T+2bIXj/RB7hB3msgLA1nSkqHJG/qvXLCH2RP5MQApYZ0K/xQBMIfLY0DlEEEeiXgkNMcUBO
OkNvfhsilvBZQFxpLAJgilzYCtg3xL+OLJVbldSVz7vfK6kGze3TOAblChU2DsoARJuKVWPniEcb
QeyPbQZW4XrrVsAC4ab9HVSeRJ3wQ947mUVGkAZe6f2emRa6JnsaGZng3d1LD71TExwd+iKBBQUN
oC9bY1ViC+c/Sh8PCwWXWaTTW3vkdKNzP+j9a3byn5EiCztF2juVBasCzdh5wfmBnDBcXmAr2Y8H
XULGclyYfb0HYi4BYfnT7QMNtxPxNwIGLcXi773HbjzrgT4nFckEk7Bv5+JraYk02Te0sKhk+fSF
7Wzw/bdcrgwGSw+gTaD25vy5F4gV9hl1CLo0IC36Uv68u+YsL2axCP1nXnCY1c1fsBBSJv0B5NtE
ZBs5km+MqaGsnS0xH4JQttXDjhGauonVSJxyaybFYY/Sgm63fbMKkd+Z/tFWDEkYd2Vtb49Sd7MF
g3G035yd1KlOLCHoXlhMV+WbkYWt8hcfOR/gSrc05S2CHlOX/kskdHOTiF/wX3bdHMmTqO07WKHd
JKeBWE2yWPwNA7Et27Kc9t8qebU2X4HanvX1UAYTGoamullNz/xzYlwUFTgYeLh2NYHFAJ714vtw
mOiqqEeJffVEjXTvHswbBiaFHBWj/dYPy1iMwvCraDgFmjeBH1WLOYlglCtCVCcdNWC7X/hgsAtt
4S/HwguHAFak42AsWOZRyc0dTfNLVhy9w+JBwTfah24xN7x/d9NxMNZq6AGCaBuwiB2PHGUbI9Zp
6oUnDchGrmNbD+EaGe76MA3XHgWMzwuO5MG9kO8t0uATDnT10YAgJ7IP1C2j/E5iE7izqm0y+DZo
yqRzE0oxeW3cWR8ygxtVKEzAZh3FAOyQruosniGNYjnehF+x+Fv018ROBKtJzz2KuI3vpE1Ort64
xX85zF2gRMMpW/V+Xo61QBcyvWMAUoKImL17U8Tj+tHgIVAfMX5izcc+micmiDmbzFIKSitV3xS4
5nul2JO9jbld2KCxvLQROiQfbII4jZtitJX7RwPuMF65qzw7wezjWQ2YaiC7mwUCOiUPKXLjYLBW
4wAsft8H2hZuEX1/nQN+fyrKcv40TsIHquzLFYR2AfU0XPpH3VsGtb0EyC/I/x25yTKeFEd4lxPk
mr5zfcsSyP8rwYfoXp9QPN+V26AYYmZ/Y0hgU56q0wz/5wxJPvICizK6CDNIOGkR0YDfcf+YzCub
CsSLp7JAjFrcnKU/5o6ya1emzKKPtGoLnJO2wf9rWOUgeAloMznPwQx64Aeh0nV6QRqO+WMyHIlG
vDh3Af0FM3VMcS4iLrsC72fL77jhF/L0gYaasQ9+rcc4L4+soJbmpqtK4MzeykOUkD9Kxi825RB9
/0OSvUFwxH17OQ0dLMfn+IORo7C8SC8EulI354EIXHFWPOXY4s49LdMYs7Kq2EXwyXqGGFUyomKy
G9HJFSxew1Jn7lEfaoon3AOZdlSV2s4/bFVGHFZmBOJTlXHpqyqGbPH0y4g1ns2SA3EZa+z5Wk+E
XyHN2abpfUpNNG3ig6e5hx5BAU/7Ui0rpopEOCF/uCNEflemtj0OYWRp07q9UVgD2wVJwxz1clTn
wRDHRPIa9ddp9J8qFm2ijwFQdOtYeOQMimxviqKzqqMsfPXLZiXqtTSxw/eiBNPjArTI8rQRRA14
wnHgnVdWA08hnjM0f49Dz6OI1EOup62agIuSItoC4SQ9geU/vsaAoQplHxTeLesZbm2mTLmgWEpx
qWk2yp47/vRcJ28fHP7B7GMGP8rnUh+2gsT8OicaHmCQtQSwGKq+59ud8vGQCy0eYuO3KYTJF6Td
MTxvppe7i17e33174r12/kZKVtBnkwolaZaqe+xJr/Zh9iOJq8LXbkeCCa9QxAWNjyITaIlG7qfX
sq3I56Dr83X28Ht6Eeb3v9dYM0PK2II+quY2DylJ9ZanxznWN5dzsEb7DfO35XNu8EmiTWw9Hkvx
854PwQ3mxr3FqdzBYTb68ACeH83wwfmUarjitihOvEUnx41IyZsLMyQ6hMxWOcpomcQuEuYkCxUt
SRXwOjba0Stxz4WIVEPb/qNDjnuRv80u6h+TLesooDIKPLT79pTanO6ZdJdkXrIDw7QRBiJ7YxeI
exteukI4FZyj9anxdm4uJ401joEAljXtNSiXOdJuCKx0d8R8ah5LJbKmvzAGRMKbro3lD26ES8Xk
fRw0l+Q2ZYnUzmcWwANuT+XJI0nZ6NJAn7/WGwKwgk7E8WAm6FVpPZax7c0rCsJVotBDuLIzf0uP
bSJWuSGPkZEQewqHoRckqoFLNy22JR+csX2rVfhFx7Y2WvOZpbQiY/b9tmDy30Te8GwmR9ewT/lE
sqjLmTWWBrTOeoI/OjUBsZNYVqKGN7I7a62XpCUru+ZN3OWcL4I0XkRrr5pJidGKhVOyWbK0po4V
DM0AxNXDlEjYkKnE1pwSFUe9pE0bKDJ9hHi0yWxXh4pSddOPSAOLx5XOfW98yEfQ4uRuRKF+1W/7
L+0ZFK8HsRGFdC1QyBmqnZlB08ajcf5nzwwQgxhUiwMWpqVXzEKOUGX6CIVf2INjAaJozxj5Ha3F
Bi2r1QKtr0LA66H+7WlDoEoYpE51yQFyCq4mUb01YIH3lrES9wK8dcZYm7/uS1OP3WwvRSaNFkR4
I1ydjQlgPgRPqI2EGuO3nyUur6jfYaH2KWuq5cJWLSzFr18upPguR4b51J/5TpzW2mc0wIWEh8m1
3bEsM5q2SMh0bUk5hRAqyG3/Aw8ujY/UI/hhUCvIy10gXRli9KH7sHdABziS4E668OtnRu91vPpH
jFseh/9ortluH9hX1s0SSYhTS0UkjfPZvEP4JXirnSYkZ0wAqGqZYhWmJhtKlogK+DErZ2DjqfDy
KdQDB4u2dsAWKX+mag0UaTptncn+PZ4Bhy3KxUOKUVUxkL4cFHtdqk0rS9Y05VNx5RJdsA2sO/3y
zlnmAaFovUSW2KZSR+7QJlBDjRqtttqlt4Beyxj/FMJ0lqHOz/yUJUPzzYTm99a4Oo3nsy6Yu9TC
YGZMYxN1Iaz/fxv3n6rLJvWykIF7wXGxSR9K9X0VQL51xo3wE+NWrJIXzAPbvj5iDcvidBwv4H90
I/vqdPAWDUM6d7OsJ7apNR8uu9sh6n6rdnbXZzS9iJmuBL6rxAxEqWw9bYyw4o2hY/ujjcYAZW2y
y5/0Fa2usydLduvA7NhJjjfRsf8koRXrxSDbrMwYdg/EUiNeshnoKhcweA4RWQOyLfH9dgH8qqH/
x23ei0U65mNsoba0xbfYSP48U522eCUsnFXCQGshe08Z6o3nMvaE9ctUxqn376PCs8gTerAZouFz
KaSX/42CBx6AqiKMJWYsLrdzifDwCGE+DJzk/Nzxi5d2GPRzJ4oBehX3s7c5qrfLy9fO9GAmHCN9
P9w+KbLzXur4r2Kf/7EHtINqEw8T3C8q15lUhpjlbIsm2HaU5mI1ZaZqOEhO2Jz1CiVapCxzv3uM
l+y8wfyxekJlgK4+7mVl9bbCwIFdEAmIq1pRNeqDJZ5wgmER4x9NjKt3jgVrg0CVTPDxJWefg3T1
FtNO7SEILMQfK3e9iZ3sYolCiSb9tiLdP0zOrb1HHbLjJsarWAa2ADOrpV3EyQ9mmo0pgfq+nmUr
O8U31REFwe9o4tHeuMkoWHtYGj0HnMUJ27R9Y3XI3YvDPwsYTQvR9IXf7nvljn5/xN6sOy6iecHH
Jpr0dntdo055rr9WFDlEm0liv68E7pXfDHZt030uEwCKijHfEeSILXJcWmQHuIJMmJqLLicjNHok
Mn1b3UwJ1zP5BtLVQ+eChOMSVX+NBLhnnMQnuGtRos0gllgu66S59CsDtSeIXqvSJx5b3Dsw7X0F
Xb87ey+66qjHSIhC4cwe7gNquvPw2I6iQJVnkGkEDHOLiaRZR7v+AJ5fOdblcd/W3m2xlSda+9DF
E2cpzcEJv/GdYryJ8OeF0Bw1/rPOmPCeJtMBPj+ANyYWHgOPaVz6+ElE6VURc7CtN/fj31XIx29G
WS1wKexmfHtymGc7MOzXNZGUmVJ228bRbZrMAXxWI9/IB6/P3PqwjU/Zt+bEFn/tLED6WEQyz64u
FxGtsbtx4PnsAO/NTa3O5Umbau3wul35N5lYylaJtb7pLqupbd8Y8dBdOHOvZB9txrfKKioEsy36
q5/qHTn8xXxtGMeis8n0ot8ioAYzST3o/iZJBy4/iRS08JUKGyAn3YBNpET/DYX4NvUpa3hYsmn5
8Y0cK0KsJpLl6NaCVICL2Iw3N5+wdDwXrqXwSl0BACtrnmbB8ntzddDZjUCSPhhvPZTKsFIPLgGA
7URTZl1Gs87trNf9v3Kr8vypij2SzLAfHgfFt6BOo1kKcCQrwqJWp7o5art/VZn2nxjqKx2rU5yE
Ht8MImCChupDy32PPxBpAe1y++DVG9qbMiWrU237QKOu6gjKSEJ9t/ugZZEWpwKJSoUb+WgbPnwD
3E9Ehbuj26hB2O329AjkGw93WBX3Wg7O7uTyCtcdvsB1cj+0gFVUi8M44JCUnaJ7XyyeOkhVZQcK
E9wWfbdLMyZ1OHWjVKdk9WvDYcturVoIPtbtQlMnIXGLdVmieZ6UCrbh6r2fTLCYzdkFHzbLbQjq
ituzVcjNN7b7ij59fZR40CMvQdxwX38yF1ogFELlvXY9E/Pm8uC+/i6toYXr23KntGtXqGC83SHy
QU4IzlkOuPMQRvqZ7jb5ed22nyEDQCtk7hGmqeOiSPd/8c61CwviVIUfTjdv95mf809/qv1VxMfH
YWPniWwwc5d/qeD8L4p3ev2BI3lVEflhhTIvCvKH9HXm8sTaImnBdQhSgtDOifMTxMTxmTkuvlnw
km5ctZVn5JVln/HbTNwehYvC0WaRO4DCfgOMBOyMIasQlEnY5+AKYehb4/f4kG+opfUEG2LDftNe
NzYvQKhP0jCRs/0YwKcpvJZ73iM6YSwkF1/CDCi3Fc+1ZlnYXD4amOQoc0hRpDZ616m+nsEETys9
+3O/AHmbWs4meekR8oXVCVxFd1zcVEr2O+dh52YssSXPOZbcD7fZmksqIvdGgD5ewdvNdq8uBOXU
N5mcxal4oit4SP6uwV4VBla1baLvpxeBv9Pc9rcED4f0SVV/zzIuO5Vmo1vjik0vWt57i79qVrVb
fqnLvRBcdlXKTCCtnmYLS2h45oHh5Ck62FpZ+tzxvXp8fmCKJO5Ubp9y/DMSth768T+BLBrvPZ/+
rZPYSFMD7NXj53JP590dSmL/Wr97prGUyzNuR9g9f+PClwKVvV9rPo/1pRkcyKoH9dkF47h2gBKl
t3nPCilKAm1HyUipV7vc1sTSCDs5fAIiomr2i6OdI3st8krzlb/t+RepiqiXE/atiDjaV2y+HgVm
UySlx56R5rhnunOR+EsH/9uLqkya5xEC9SSKrgnK8twcJ6IrAs98K2JEIzZnLoNIimppCSMW8n9P
qIo5WrANVqXzmm1QJFralAAc0PEnLX9SHcpiWWF9DvSf22dTQe2AEDoknmbSxs57ZgqOMpL8xksw
rqFststbxXjY6EGcT5ARgeknbGQVyf1N3KrsWSlOOU9/anF1rtJPAXpaoISTRHXNZWZPn0N23woK
GdJ6dd4TRTEqaFr/AHlMX1bW3QHhG6XAhTif4l/Er9eDaSGnydf9I7o5d0+yKf1aZ5BNvIudAq2E
e4nocukF+EahrkOZZlz2UQk/r+v9H1yTgnJJCDZigYlnjyYIrVozRD/wEztfnWDbsPO2homZae75
IIPm3ieHGq8J/l7TXVVvfYaYYenidzHGXzhJ76tDCeyIY5m7mtUFAY3qMJWG/lmqpG6d0YgF/MB9
eSiOJFv7TMO3TfdHT/qnV5X0FXhvu4JAq/x4MHkkfDHele/v7KuaDXjzRoTLQmy81DGO2eiBQYzu
qmXFVFn7Wg542q3PtEKzM8lZBWelltrlUaYso3+00OEv7btX8hV5JNh3fKW4GFo2k+gUtC4M7Jpy
jiQwDIaby+faoG1w7kdMDOGPGlo4j3Pv0iICeXOqvFlbphW18lETDgjWiqbyEZpv8Jpx+XfC+9nH
6Z3xEYhaxjgg/NxYONP1zI5b1Nf7MhJfyt0PI9clcbUrxHpY1GSPu40bagWXzmBpJ+l/ljhhGHp6
mSNFZQ3anSpTF1EXG8oDB31ZV6P21qWL6e32/tdtwqhF15hv1LpwzZRfd/CX4QdT8dB57a0nuEG0
G8MkowOdWvdVN5o7hBiiaTcTRbLIaDAdbp4DAErWkGgMfN92QQzqMre6y8QTCUL5LF1MxH0kSw/z
OnkAxZrOWAoZsa1lLTbrJj/GXRuIrRAwolF4BuZTHsiH9G4yZnp1X2ENKijZy9Vhu4qXQVsh1nP9
GP1UHvc5vKipnZlmYLk7ogCREjyOqBsWt7VRFBQlZDADQXa82kCJ6X7KhwURkbZ5VSTJCZlsbkG6
CrGW7HFKbBzBx3N6X7ljEsxZa0CUYcjnm90nD6BIZjD29+/jNUJIVBYDbMrUjaPjd2pQFrgmDxUX
c2DgX1xnaGWMze1ys26xcIX8xqlBiJPZw8mugd4y90m8yjRvWsmojToHUPYjwXW1V4SMYKC1c2Bv
iYApV6qMVXeDouCCiy5E33FQgIa7eV5iRTiixB+OqP2lQ2mhXuVnFla+RsZk3wJdgv9QUWYOnoIc
8gMQ1KK+PmgFKEjSyHe3MHOJ97d7T+Zd94a2MvOY/JmA9RcmPonrdRSSxWCK9czEkKuccig+fi27
GGCbUs2EU8mkL0STORruKsuQAlv9UCOJ3n7l4HOy9BMmMv2T/PL6ICdQ3XetE9XMkX5Aya7Bp+0i
h0F8hR1vjnI5ozDwwFMe3HCDYhkhDnzmZb2RvjZOBF4CMUCnxSOaOY9rD6+d+eDnIsIMXIA7pB4B
g4c1ttarsScTEADHRp10uGdSustJyZX49bvUNyapxPSBumHuS7nMJZIFJJ5bipK+gEjwYM3pdgZh
XBQsrKDPBXalYwEnFQRQzibXlnztLp2kX4p+7z1TXoOZHyfAuo+VUG3XqZS4T9r5EGGRspCotwo0
0QDZIfiTLvFw02UxeygsYCy2987/ox7LJox9Eh0UR4bSWjJlRhrLfcd7/xsZwwsIXE9LNK/tJQ8B
I1tUO1Dp8T+sfPNPeukIqwehbfNeX5VqLNUvcm0c+rmSj62n7Fo+pnet3GRPaM0xO7gNGyelLJFu
bAeqzdZqw4C6JZJQg5UbDjRSj0fp1/T6xUUHxipSzxwM6/mrcUtDoLcTqYwWWoQamXRCwLyhy8PG
YC7E61sOD7QiVy3TnazqkqDIrBBWxDV7ofefHbYR6kLYGI92zvSRJGxuLn+Yif06wPICd6/ATq98
Bw4xdiEbg3EfvobljR8MqhriwQFDa5yLy0TGxLEEDya/E84DaYAmXXfWobQEAw9YEXJb0FkXZtyB
fPr2q/g8iZtyrTGkTYbxo+bLqtVnYYsuOLTVMVN8pEr+fuWDJ6HZCcYvBtZGd74ZWwmhU3Nz8Jee
5GEPHSvuN2N8aoiQR3ahOqh1Sh1ZXNg5XhgVyEw4QeHC4PZVLI+lwVG2A5j4W10jB4S8uSPvloxT
7VjFw4ogEniwBhGh7iGr3fvFRfRLFNEW0zbo5FBYzspiYzJYpCAmwlxdf/bLWD7vskSTyoyqjJiw
CVbzDs+3Px5LFw5KWuerJQ6oGg60bIVDU9si/zswEzoyQR8Aa6YACqZzAv0LYGKYh+L1a3rVkvu6
eVlK5AqE2Ac+KZNp66KjXOclw3WdVpDFPcaXDLV9pjnakPP/Xrui5huhxH/LKX/8toFoO976azwN
dSq3WGtcYHzEo/HEs9qUGcAB6YM66M2Lp0KHM2wDU+FS6XozxQ1bJlSnRKDWE7fSPR2L2wZQQxyh
VkNLLuRKhlsPk+JUaj1PLTLZ28+rgyARsFZddSFfxOLVDsfvM6qPFZ4V3INWqzlYELL3RQfFjiQq
V/9F8x2IV250Ux97o28K1RUd0MpkV7C0OfVu11zLVr9eUxxdr3pvo9zN2xULGEgGs9Mlxlxg+eaC
WU5MQ65n2Erb0/DdMBIjsDM6qeEr+5NOJEnioXD6I2XOQa4+6o/28BaU0G+RKRCgmhzM5CV3aW36
FIkfSSO2pUdPPPWT7MB3ukkb+IKvxg6P2tFET4G9NT4qeuOi75DoMM6ypzWNyelm7kuTU0RqzpV+
dGEnwrOH6s5UPX5WRJQNRrnBDeUFkBHRVT0aCSWl2YDkPvg/nL0k3Ha6FrMwyQntukOBTLqSjBD6
f/4xlT6SuxwzBl7fZuydfUubagrlgg0ohREgdp0jpJSAl6j3qpS3AmjVx7N1xB6GkjpIIl31Ktj0
m0+O1RPsEcXI3laKj96FwMwBGnFpzFCYPJgH5D1RmzqPrK0Dr9W1SC3O9oJHl6qWcj2VwlfbJuzX
+3VxnN4MmIDM5wcTPn7eaSOIYoNkWSxZO/t3BbjVhSHma+Ujo4gTob9z2U9JRM4TsOx2/3jlL5e9
+IkTH1GlXIUHJEkrpYKVC+i48jpgDIbNZ50Y0yPMIHpgsS7krsDBkFmdGvJOSL2pYZuasLN6Wuyw
C/WV6l6Zyujqp3+Ie0poFSfUhsnrOx9vElsJqeUek7y8QHWZB13l2PQ1OUpxx1EKvoENxhvESXBS
Eb0KoRZTNbkCQ5/nt4SmO3c3DjVpWdQsX8kkQP2FrEFM6UCs9A+LU73UiozO4sYZTCUFPYU16o7u
YxXsDLHor1/TTAfwOcjqM/TD9Huz26hpw8O/iM3lzTp6NYnSRrCf/uA+tu31HPzpg+RdemuBm+dV
zuyLVhcMBhE7NRW65aAvSxoI7TggSXHGdJJwMIC3+2lKqeNmSKVht0A1aQ9KsmCXxJP2evVqWgFZ
oJ/ftK7v3RDb3Jvqi8bLWVUZDRZ//rb6fYMpXBiu2c/nsR+vbJiXSC20pNWDZGWvRmgNqINQ4e3F
3s2BPnM1RM8E0IoVN06gP7Wp9urNdV8M0ApfLawrlmXlZSheEPJlXHOGddqMiRCPDEb3lfx+doiQ
/w7Q/pzm+oygB6dOxK8VFICtjaHdwBqlfrxMV7cCoLWXHd2R2BtgQRGg1+EZUaaAukpkBsB5lsNo
4szkyvYDHAZd0Rqzw/+90So7mdtKcca4Oj7FiM7BJay/xJ0CfzC+CpBzhH/8vwSzowZ7cZqMKHec
qc2pcAJ+/mvP1F/U4PsnlqVsDK1abE6dE1Iw1FpPJMjDjy/t4sfySE30aAs4YwL44Qg/vnJ108M8
7ITBA55pMKaR8KodEn65DQPu7nrdVIe8yksEcGuRlUAnCGFwcCLOST2LLgbs5mFCflXTi2c2MLsI
GzHHjjtWF8EjrfsnPiyxCTxjAlFu1VXX5CI5z8HIpXzXjodeOgPfAZOl+5/7lrilGwhmu302+NXH
D/dChO3jPhGezHS31/SCfuvXPWdNCe6qNnUqkJtGjIURcxXRMQ13Uaph4vQ77fzIX+Ng96caD+yl
VGBId/EYEESIcNbCWj3ASlWBZM32DZi5XoZFJxAScT40ku1Gh49wTj1WYNl7vk3mevtj+YAndvh9
8PgWT3h/Qv4IToZiZLLzjWtLqNHe6sED0rq61L41YvkNrLyOBCBsrbs2ucq+df0DXG2JeQ4vEEW3
GFkC4jXjGXYXnOaBMw4qii8gvBy5QhH6/2OMP9NslXyvA+knPdbUS9kDnlyFAig5h2o23drXAsnj
8bKY58pT20MrcUVwalvc4vWI2M/2zH47Y5dSVgT+6ZMFnZ4t04djmqh77THAoa9X4mIMaVgva1i+
5dJB0Nlj4SfdUl1zt0aQk6AFNWS3Q+35bxmgzSHECQweiXBQCbsCtSA7JC/unMj1JITN22YCKeqb
og9HfrzWHbgL2GQA9DhTjwXWTxqnuVNZvTXBY7IyJL5PV0L+k0Us/3q5qLTmA/+bMP9nP3aC/Oc1
L2qQG++uv/PzjVki+cVL/1plB0XsMgosl1pbHbKt8rl4J14GPMD0ympECamhbzo8WUutGnUm+rSJ
GMUn2q+/8dR8oRQZt9TXKseI9O6yI5wl48C7IlDr/zmmk+2HBYrqt1QhH00MfxQ2270uYB9BagoK
WDNZ3sha0nmpxlqKzcZ0H3dg/yDsJiQOET/UTR11Q9KOjUYdsD+5TSBtrZ3xg2YfgUdHtCTQ+9m4
iy0odsb4897PQnkd3r9h0ytIPI68NOSeymaLCM7MTMGz9uJ5L0AXvKh7S75Zc8mUPg34xZk12fGj
GshtlYsK6ABNU2O9A6FtzlfUlj93Uusow8lBQWZfl0zgXvvEDBq/hOyWBXP2j11F2ZpYzvIs0wrD
btVoSoCzN3TOTAmERROhpMb3XKlKCXdxzOkWhhB9Fr6SqZAvPBlCqKzB+0OGwehDNubq18dCmyC4
zTIDPuc8E47DOu39HHQj8MHsI6zkzdtfsY78gJWeGDxC6SGY9qvzP4BudMHqcaTBS+A4lkxSgBJZ
YrlW7pfFUQu1xJzwc0ljZMnAQ9P11V1FqddVBBrC0mMusH8y6qRdpCv4GZYc4WnLutxlgOC7bTul
Wk65g9QFdM7lsAepj9ugxKfGXWiaA6AuC6Ct7h6e5z6GAUFH0iFRxX53d2ntYf5IzhVzY18BfspU
7iy4lVFNzzy6utzYh2V0WKBdE/fO8bVpPyVmYsK6BfedD3BV0iB+jqEysPRs6gMqd7Su561lH8zd
DH64HH25+O/gWLDTO1mv2OU5ldmZHhY46YdgVyQWYxhrkdDNuEw1v8w8YO2SuouUPCRUmF8+RqoC
XvbcZIpMpP1Ma2HhMmKfwUbh8AER0xDyIj6Y60gZ67D1zikYK18Qr7k8MXRVDZ2/Dg02pqdI6dij
U0l/dbmp9BRGqcBS/teOa+NDR2sET075FQ2Trkom1wSjjSswAhrX8t7eKxkez+sqGRTrbp7iZYNu
qKjbczWoAXu/ua0tw7LKBihOITxgzFH+Q0+9WxcSMVI2MtJbkzd26SDtjioWsGLNY7cSjSKTJnGR
m+pHKLBz0NuVtEJVqaRliQZ20A5JxHnzgtcHJ8KScPFPbVThx42whKz/dPD31+fdlMTPRllwlcIL
2abVaUM8AXGIv6NHnWnRkyqiiRoP2lUOa8Px//UcfKYq3XihVXcJ0jI6TzAT/f3DDEqi3Q7RKniA
XQgjFqgVMkbi/ciqbOjwdIRyldqFl8T5+YpmpboW2N20CU7r2fvptqGe5vqtcJHS7nGgzpHSMDoY
0CV2af2IWR9C79IBoVZfFX0W7wEoAsOFjKewsZ+Ka7HFxnpySYV1878m7WMvCiLiplnR+yYs/f+v
buEv+FxJxn+sQguNu223tyOT3o7I6FN8cHx8MD1HKN6PN8wshGGhCWl3VbkhGAOFDJdieCekkpWy
xsq3beJTNqfjG+78UkUKsBETL9akx2Xe0213Sk4lY12daEWr+4n2tlTzHe85nwHMnYlGmxs246gJ
VDPbLQHrKJjZv1WQnwL+liVP6Ou+xWKlrjgjMAqMU/HzI0DBf0nYo9i/wqC0ymAqXA6FZGPJdhpf
/UYCRRuKR+8fQluTHKfvzSz5ODeIoGCYMI3Ce68vK5yE5RN8gJxG2zx9VFJmGUdBSWlr+vO/bgwC
IhyFp3RnlrR5BxEhmvhGO75v1F2ZFz5imXWpnigwySzACg5sgQWdImSmfh7Mo8g4NfuYDdRDQ8l+
uodG/3p5nJvRhUNVou9gdQWHIQLigrgzNSsMjxcU697naY9mCNBRgr9HNKIims7fU9HEyoJ6Yr+j
btnzi+PhilYLpuvVNQK4qS+btZIpefD/O1/CqTFA5Fh3VZksw6khPxmfbDqVYNaLmUxDUbClETEP
qoil2iFu4AMDBP3/sslypqZvghmu8/jKb8crd1p6iYVewXVL2d2tK74NR+F8iDlRFhLIWMnjADzU
zV5QlDONUqaJE5NcN37hn1Mdhvdl1iHJIY7wbZ1mUH0nJB66g9x8JOyl9yHvz1REqTUvPZbU5V4T
LZVcBij98TULCllZQo6ahkIq9PtPEcW5LMBxZ6Zb9bHalanTPGClP6ABN4oiQVGasLTOC1qUS10K
G59w70xV9S8KOJWz8oKLB8PloCAUaVqlbsT1DwgLJAl8rLaOsYJBshGk2JKU5vrbP/5f3KLN2pz/
OZGFb8nSus37TKG0ECV7biuCM8S7Xw+NPxZvDfBD8Xcvmd8JqTecACZ23PH9DRuOKkI9HWkAfycX
KgXppgk51xq7wWI2Aqtmzz9lbRaT0hHNMMvWtp/6rJCiET2KchAOMK3no1Ul3UMvOj5E9tgu0JNK
taEW/tDfAKGpNiuYfwf21dpk1WY86QlePZq0ANbK/lSIrh53CB2Dey7O/q6py7vhs5XqcYFCTXkr
y9V9ZZgm2OLmc/UnUAduwyLLK+ipynYYXhgUd4lX+R0A3eej0m6C4kysbEKl1ksCk4N3tpWZEQDh
0IUT65ih6uIgtoGepR/NeYgYO3GN8h05c+Km6aROmeWd+yCKcG3Kstir13JYV6sgTw/dhnK+gsnT
UnTwnoRA/snuzrZ6rtOu4NS85Z4f7He0/3FY+JldlCoiTG60HmKQMkEYYGZAp4fqJGeGS3CEs4LU
gayhwlJvpXdPiO0TEOnkTJ95FGpuX1YZwE14l/dN0hWMXlP5LRojk0dFRYFsn1G2KAkIFNwRu7oP
ewwk1PRXVJli/4vaQ7jXBsRBlotBy4bRYDCtyu4lLZ6zacXUrJn1Pp/7tOCklBf0uh1lg1vtkH7g
+AM/s3s/X5H62mIioRkJeSi/bXUmIKzPQckK/GQV1ku4zrTlNCwai+vgxW9lxNaY3jTvzabnWpGU
PPafRW/YU1HuLlGUtGwWzKoYslFlgAfC0nbyuBUA19pKhdFSVArCIc+luh5014ycfIg7Vzhuk+Ti
MvGMfid4QnpReZCgMEqEFaMq+9257xpsJVoNJb3BVZdrydLTQCsLDbCMQedEjdPGpq5ymgDd3aJH
cmKGNd4FRAddcCDwB80+82YyCFmnXMy5jO6gBxVNPxOLxsSafHMa/ypXcJbX2sjvIie6fbTJ5dHJ
hyj393hCDbkPKVgTB2IjHNvoIZ0yzwwOd/kQqSW8pBSQP+Bv/v2iGHJhJLs8FE9OVyo23Nwq/yZj
knHBraSCjYvI9lZDV9VIvHCj03GJiqeG3FOoW3VAwQb0VRoloBH5Q/8pIbZIQ9epUYmiR+27o5f7
C2Is00zGQLpxsD7ig/03eUWD32TFVge6rVtsFR0/Ww5a3QMHkD0H0LAFBJqE8Q2jc4pxKYF51j2I
RtXZpuR2RSDrQAbQ14Hnvp5kwu4GRc3g0r5mxckuTumlgGMusM5+wyQQ7uiMpNS5ZrMPP+q/4LHY
z1WM6W6p2H58F1FyJ/Z+hO47czcrVPYstZ2ANxwDzw0SSsp2JbqNuXUjwrMcS/tWL2/nlr3Gx6/t
s0+lrjiD8C/Hp326L6izJeD9T3s89IV7m9ceUY/YhA4fUuKvyDhF87HBhb67sHLdzh+zLVEGzRql
ne74oOsbXtIzt9YziDgYroR42YmTGW1IAPKr+Y7eKNK0eF5TfjF/jMce3Mxdxg3idDCu/Kx9dpaa
9VOF/c/vvycx1HJ5tpk3FyIbzGMV/Qgvz6z3cmBx6M49Iew+bllSquoIvkZFPJSg/NeB1pVnVnNe
RVcUsSQeVpOSOS6tKSJ7j3EGcNuRDK6D/nYATtAKRGuITQhfCnXO3X4dAly2d6M8oiHjjfAdEx+2
RRU8oH596lmOfa7zE62QWxua2dk/PymX5f/80Aq9TSXOt72ykGmPacIefma1HgZgvPXibXB9igfr
zSTCftCb0xGT1WsnybZMxKV+VjN0lIkHuQO8pOeXcYbv50BLF7356xPkBf6nAxCgviKKFJgm4ncb
iCMfiRFZ3kR3XLj7pvLIpj302IMmCym+X0XUn7l5VZMDepGnye1zWicyJ4YirR3A9m5SZgl6hbdm
i9b54kLXunkZX/9B3jmJyPRmoBWmhJBeShtH6nRCwsJ7extIET25m1vvM3A8+TwRSVYnTslc4oBa
kgEKUD1dyG7Hgoyj2eEblQz5sczZw2Z+TkeN4NKMtBZc9G9LraqqHX7roMqpGjoJNMhDCIlNbUQV
UWqif/HWioTkHhGvzZE5p2uOl8dAZPpW/L+Q2wzhjCuLie0hDCnz3glTSRlimQ/UF5HatB5ozN/c
5IGQ5nZMtCCn7eTAVJ+HS7ScGbcS7fhuXXfiVk00lkDA2jXWhk7KsGx59FQdCtZvfnZx/jPPEKdx
jWRtKHs0YbT4gRLavkYI+i3kLkmv3/jrlIOOAtJsypQLvIUSvRGtuVIQk1g9CpIOQab/pNxDgKkS
PkAO6sAWSBpBvtG2iaNXe+QoZ8vEx1ggadodS0ldqqaYaeaphWbQK6VgwaV7pMvqNORCuv2bDFMK
xYJ5RUODEeLEkiVy+Gi9RR90g32BXHyZ9Mo38/IWFwkrkqL3DKPa1euYID1aRBAcdistvzIdIx81
NAII9Tfw+QHvIdo0mbf16o7vGKxHbjSDEAFM6Vvwtp4owAIVRDdSb3g3HIEXdMotx78DCQCApMTb
18yJgmhjBeDoWqkaWJJbn0Ka08yYuPH3gQtAQMmGPXeg4PD6NPXmAtSaSLSmV0yUxRAfEqkS8sb7
N/F1cEeUnfCkoUOJH8NpeRkZwn79I/h1CZLeYpvKotj8NNcGvh6r8zmTx8AWXWtLKOTsvF8Y7Sl9
fSpnnKZmiGgH25a3B1kxEItr48pxVIF4rLsGigyvd+GL8ufIShBJyCiWTyNiEzWJdvE5q8RppO1h
xGkiEU4JAbFnZkvJndijsHz+mdG29dC44gcs8Ztl8KGzwE2vv6DGmc0wus42k9vdLKM6gpenoySJ
shLZ6swuNh79D2Xf9KnfiFyR8sdtIu3RL5iRO8RDbmG9nM/6l8tbhS9otABbgwy2Kp1F9EUan7uu
uxqr9jiMAaxE3NYAZMTCOdIfAOeIThmMhuuiFJ+PYQ0gRSgT7kNZu/mntFzxSoNNkkj7T3B5jjAZ
DmPZKWDEzuBNmJTtsfzR6jzF6SePPb9WFyrGDY2yAPXN+nu3NQbFYRfCm3+eg7ipDHctZokb/3P7
j057+OaQQ4VkuQRBYyquQdOqhU3YiWn29aVpzyKqwgsLj5B6oi3q9MC1FZfmsafeb6XFD51viewn
qi0Lwtr+yuaTPdDWDJLKXVzlanI6DMVGFOp5v2xVrp0ieRv6fvn9ZRFDvx9z2LYMZGTbLfdwc4AA
hSVlIDreWClNj5rj4GWx5eK7YNmP4vxl4jKd4DFZ7BIxPyinesR8BfVVVG+WgmR8YA13eVaztEQc
Bc3GALbXMh6QiSriT8gV51ncI+5nEJQaXcE5EBKAKahY/w9y0jgBHX8pAZJ+F+V+a+FVx5tVLOAt
xKm8FjHjpx3PjABakQ8LlTUURFkv35iSOyiU1mgZrcPMlYw4f7tbVWzAMg6zXLo+edj+K/a69F8v
1iSm9FLjKntsUb55mRLZD/Uq+o/5/pjy9KSMgTcCmtNfT6F4hxBrhDQLB8kf8Bmki44kdYWlYIYQ
xCx1lScblQbwJC8HSuMxnMPO3jEZR1DmrQjHda5tew//JICCMWHvTErU0ePT5V06zajX7CwNBWev
UewrKo+xY4ddW+7noNMttyBNnoAKQdlHxkCLe4dCoDpbhn8m/ddPk5aVEmeVaYlzDad1P2PfZiII
b8mhocc+DAWpkuGNJhTSSgNtkJ32VJXmsT6D1wX24Pi1vqZzuhnNbLPWxvOmipBIevVKbdCYd7hY
8K7E996q98VDSd7HLuvKDAEn7upJKIbx8i0XB9UlV1zmihCDKzIAE+NxL293/oY5tclSwQgIG3WB
PLxqPscP/9mgI4heA2KDb+b9X3ompEoiTZTz7DCWTysLRTLAlG63yvtf6gilKnte8uG5gR2voRn2
T62EIbvnFAZaFbkFRHESVCIYycLQufcIpRvXeezBFAnyVf4ShezU63sFME6mXYpK7kCeo1yZcNiP
rOAmHpTDBVkvwXm2oPdXe9gvv4RkUDnOcWSkLG3FYlRO28Tkp+IAL7r9zBDVXN4Pt7ilS/cst90r
wt/tbJ83+Bvb5blw7LiJylBbAwk+D5G+D+ZssTG4H5HaCfFbKldvircvMk8oUbt7XNuCuTl878yq
QdNHlTBbA7kYYqpwgyUSlgBGyIBX+mMlplIw4fOWsj/x/hpjB7twPB3AEDOyzQgZoo4kfYRcG7Up
T5eW6bjyLWbYEL+s7bBLaxjTXde/ZDMWtEcsMmIS/L7+s/qRLjLXKgxQPG0uXlUUYiDJ2c2HA/ui
iHliP/rXvrKC50v/qGDxrbPLmwMssDZGUAuqLmT2237uY0TU8Iy9rdD8kYLg6QmAb4WQawJncQs8
jvScxFypO9l+IclGAgCew0lw9BKCknD5Xsl/5gUOCON8EvOmDvZqborKTWWmMlwDnUh8ntb74SpB
xTevEpi0SstpdjCU7gESaVCSAlOMODLsAaYJ06ld7nYVTjnl2105SG5Z1h5MIHlGdwswIaKtCDiX
XBt1Hf9SRrCj794+BKTa5U27FkFUZwm0u26bshc0GgdWT1HiHU3ZKW04H2ePm2h9/eEl18UnBx3Y
73tjhw/cjy6a+A+80mIz544dPH02O2wliz1SBvYY584QftNKQ9lNV8ca5O9vX9FzJzOCsnAT+KKS
h1rF/q3nq0YVjA+3DcmPZM2frQbMsryxgy7XiX7hlNzM7124tp1sbcAvVO3xeLkshovSqT53Iok4
iRNA6ruRyb5aRN79FrfwchXJVAnuvJkk6HHLv/xZIl7AmRTZizq4ldIuxLmSHriW54ahBIFOZ2tZ
Zyokfc6hBXpRMAL6+9nVmdff8Z3y32qOR8HdQoAy72+8ftJ5peo4cIDqkf0StyHKOuJDuiKQt+PZ
mGZixV4pNxG8wN3YIRliNKbxUHSgknw/lRGHgjTo9OzClOFeTb/99JC+pvYzB6a9egvon8+II1DK
XK3WQU3EgxR+FqdKBGIDrNU8YnAfLFP5H+ZLqYzicvUZdE01Dp5w7Du2Vwo58uHgTv5yUIKdZT3c
AGSTNvsGapelclgkCMeY+EVZ3/KcoPR6rowVyyGq4+dUs5EKDR86/lq1JheCTOa/O0KP7r3yuzFy
48aD3tiYEGVz/eMTV9TT7I5p3BgReVZBjmgVfngBYBgiw62cu2fRlt2gxOHvFgiq+qfaiL+vuduY
VHSC+t95c5h6EJmiYamswRAFUsjUvcG3hva67WOkMOLp9sQZYcrAcmq5dAnFrEgsxHvcxAjftjEZ
0dRin/iA52vM2R/gI6BJUfqyfUKdo3+mRtTw+DtsKLa7mj3uVRF3W8rs8CDzK+4YpM7gbSJhZDFN
XfY0bOZgc4avqR1SdBZEVfuDrmJLCf+vY6s5plrbH8qPRAky247/Nzx9NrdRmDbv7rCzFXZBaMyj
wU1UpvmxCcCrvieYQXkAu/jGhl2/G1t5lrh11K2bb1RbrWmOalD/RR4Zs5iKfsenXBHK2xFmprpc
2zBIhG3kC+XwpR6dNjHPzYGKdk0J20ephW+PtlniRfeA5bjxDcjHFqM7PK6imPnHgsY0PWgqAoEG
EH4VM07h00/0CmS1+BN0FREJPOFTAHc28dfiGZxVw4Crh4XXAxXkV7ZZOF+KrxO0XVxjMqhYiY2L
Ee29+8eereI8Bg+SGNS7e76/ooYcBn9S1oGaoWVGzsmEzOoFr05XP+5i8TN5HKWRu6i9eLJb2390
BT8RaZYnBV/h563EyQoBhQrg4cRJhOJjvTBPTNi67Om9GBERk9Y7OgmmfkSTJs+uz74AoWIxeQJ/
BrQrd5lw4wGZfD0egwwth7skFDGm23cHkkppmBjgCUvb81r+BZIuDdA34yQWf3wRS8DdWvOgWgoh
Z7Lekp+KdNQ20fNmzII7HuhGs0u//buGJLqTxOWEisIR9gggl+v56yc7ZR9gBPt3S8yH81PGkpgs
GSBSx+BeLTGFMtDFXMb2eKsEBQVWKSzx7uTkxVL+hGBlrUEXNdY9R/6yns6u/SWHeYcS9e+ccUZl
L3labsnKrgZ+UJsntCdiDSyR++QWSD8bw69W0rU8yHaz/rslQbe4eeti85lWCyds8+e0iL8FakXG
agLsRk/sZ20jiBooW4zQE+9Oa91G4+HlQf48wLU3OPuo/pGiWBkvp5sH+TvwHyR1hjgPi1VKuhkO
/4IdsDKoNcQ81x1/rGV6fqqiCcATQfnYd8W2Z5NxqaHpSeBMwnQbV9pTdvyIiI8zq7nYQ6E5Iuqv
WN4tdinKCso9FVh5gnIttwujdlAlFZps9H2AOaWITc7pyIfXI2X/HTFpNd3DV8qAS0J0OXT4qXXm
G9PeHAkGOReMFOygTn88B2TIsHQP4zNSmCV+iXViyyuVVHgCh0dk2xW3kqgHKzUveTsq69n+eU8Z
PY52XwKfzuZWuoS/Y8Vj0lTm2emIP/GPFWGg++Yl9pAv6g4pE6EOGitKFqOSS/U9l5kE0mdQNUJZ
uBR12a0Zife+yE+3+XlPUnGs3LUNmEH2zZw7r+P/nqJapclGcw1ufyxb6YAv5jtDjC1H5AYHBiyw
v/EU4pqW+2jCWd1XK5DA437uppsXcEhTyOyOzcu1zw2ZQofeG0fPMXOvIFPL/ZhK8O0pxlQ905K+
uc6D+4kEHJ4TKO2lbu9bJCok9CRtZ16D/9B/LvXx7+tvkYKgqlOncMn8T4+TG8l0R5UdZ0BCN66R
tiFs8agTF/fyf1erNyLM0fB2YwGbM+IuERau8BWUffOEALY6jxRoqtG2WU1yM8cROTGfk57mfESX
Z2lVo2+ltMsCTNlO2SIvW21t+HAmcUjTypvrdHGJniIdCl2tWCBwvf1eIqSv/TPLKKtrtkIt7b8b
gkoOghid8hQFyNh3Rr9JpA6yg9WiqLScR23FCD5jgnn97erx+2bEULdrPsou5VUaht4Nx8u+m4yC
+61zSJf6X6m5QQ3I0csDYCoXb0MvMySwXBl011pkS/1JB0oGQpOGO8bgmvW5MZwouc3lEpkzOZ0z
gCRbQRmoGp5/x/lX6KhIwA50byzo9b8U8igZknautikA/kS9c0NGOhJVaSB5S2/cvRynAusS3p0a
YMDvNKgyCDh8VR4svSDzoi/G1XJtJXv8GTo24hn/46SFVM8Rl7fq6ZULPyi+LVVRRXYJ2w5mgkkH
qdXnoCQBO8ObDDACO09FPSUWBpV57244Iot64SUNULmq/vEepj4EP1auIKT7GECedPYVKWN2pFnF
8g12uFw5tpHRrN2scy71FaUvUzWkI5CJaaXjYIIzcxelOnCKx46vZ9RCOXlazRdajSSmvcDutOqq
mD56idaevi23kKPgVYQDcHxKLak7r3s4TcZPTltPfLOGDE2p4gpqZb8MsvKY8kdViYFZH9zr+qEA
SqPMA0oFDmM5QdZMua5aiJFg4WpNB1WkqUq1YApBsgghEcbUZTNTlZsqQASFXb+34QrFSZsPo0uM
uWCfYHZ9FPDLzuFQez7J5E4VG865guEqKTJGkIDpE8q3w1aJsnCH5we6PvKWiIfn1W4Tth9c2gw7
LEFw8At7LRM+D/w+Qrnj6HZkubs6S/unPBe2ACuRHLVWrPkXBcwA+Kqu5wJI+I6DlpG/Bbk80Qek
NmzSyUSmVnxLZ4pldTFmgwRCubfXNwGEIb6AmtcWyBQPpOOguDk0i+/lK2x71/h3Pwe7rcjnFyy2
v/iuCV+znn15E5Fg+bpkhsiQZ8nMNl4q9o5y6VbgamGRQMO+xi9LldsMdcbawfRvLtfQUqyyzlRx
fiB/Nbx2UWyr1Qgx8thMOTe4cTIJxAs15+gwUSUEcjtPdRW0G8UecAeT0QJGj1QvH19ENj+gg5tA
+yV5HV5kuJjcWW+gMlnFHo7X3oteIkjZuR72yw+b8lPEg5e48XFHzHUPk52bGja3qUb8UBoOn9nE
E5iTKc31iYuDO6cpOLJUjSsd+JIL/Ol+dHHOTYtNnQvcpk507uODzI+ciT39SHEoCRe8A+FqOfj6
Mj9aiK8xGyXjOc5K6FS/xrf0nlv3unmX0+Aa1t9RcHTJhSxHAx6S+bii0XoMY135j93ebSUoOR5T
8R86ZFxCUtQvoNpnuYvvAc8ecndp8ODPL13lKp2XXLdAQPtuyjpY5nfyIZCPRrk0DH0yUKALCK19
YlVErkcmHhgrR9AnVRUR5UDU8XgTbiL7GJW7zdFIQztJMwZcX9r5pA2K4n7fqM8nMo/yGlgZHd6g
ATZF/ovKuq2mxdJf0BI/Ihljz1cwOJdwJfbT7JKYBB8r3rfdC8rUR1n3czwks1nBowVPwkahcLrT
wRboyF5cWkKqzAPRTUCZ2x+jvZNb4Tn7rUMm3zEjmrClM5jsckdUvNf8QEHNG0GvzOERnpAZAD5N
KehfZmoMaND7Qi7Xs5R9Tk5ZAyZ2gcX5wWGjEbXdrqrH/gFEKTrzJ9d8U1mfAltFnFJBYViTMOQ/
xQZVttxA7ZgVIf/Sy5Pr0dWkrWH+5j+xK5FLTThU3FjS/45OHgebNIQNt3Rfy324DP30q8DZ6rWz
WyIf/0i5c4fjTB7QjE+FRD3b+uycvJPVteSzKsO9Vl+6172DSTfzKNqmeLcXBlEDK29Aa/jNeTAo
42Z5RPXkOc47JBNOr2OLcBgZCt6dvydB8QLSYLMmQO0cDqPKSb9ONEJUKFjKRvvZCoBgCfjov4Q9
qojPuR+IhE0w0RHye8cUuDCoSvqv598BjeJy3/DlCwJ7nD7Z0PNGZceSrW/aHdnlIamR1HiZoMhR
VyBido6ttI79FIoS6ILI74i1pZzXWAAa5ZnxRkDrEme28CXgdnhfaaFKcQ2LbjK9/Hsc42bIW3G5
/J8SUfrSYjuixAyohM1Yv6j+N2vU9MYLFBywW1vi5RNpP8HfnupVgTxP3Fcamlk4P5hC6dD9qgqE
7vsK2YZEytIMT1nUx2vDnE2oyk/M44DkF5HHKEEm7bwSvIc5UVZXsBCXXIHUxkddxCMvDPLXbPK9
LSL0lDCoUUgh+VXxb2GpcElj6/xUaZFo644lSVkLlHpP5ZAoAxVkcI93NUOcuCEIArycDZKP4Zit
cUnLzoKC0fFhF4GVjY3dsG3OASjHjoUVXvUVD03NxaUt3Ap24PgbgBAkvwq3+Z3T+p39hoHCUIeL
C50602fOG9q9kIjzkegQCMNlD/lrdwC4crge6tYfJMP9XIWbzN6plJO4UYQQ4resqYcV0gOzSrY4
q47yXd/R/0uOHzbUKkOdxlzniURzq+apQQr5UQLKD2Q9F3eXhT0Ftmxmc1RYU95pfnTXNRJyuLq4
38NqVNUfgJyKAbUJHm2HhQspVL3pOjIPyKXPG18rnzoBMRXrApCJxJO7TrR+53XHb+1rrwubin3N
1tyjfKGj72EgUQBiN26nO+c3LuMC3TwMk0QhcCaFamm4oprgHmDZJEW7tqn14zlMODgZCx0sjOh/
PqP38vbEmrQ8d0cxfrEKnFj5e2nKNilAN57oNC6xJLwXZrelUYpcYLAnE5Gf789pS58PUvX8XXVi
EVNe+fGs/TgBDwE5dzvixmxYnCeYoDPsbI+fjzTs5n1+zRuiSvMZA6PUvoUa5jqa3zDCMzGBrFqg
8HOuoT+bEhAJ3tGQuP1gOOWP5n96pNd4L8/zkNL1Lt6SU7A6UG4lxDsB9fk+MjFRV+x0DOYIWEh/
XYD5Dcuj3spYRih1fT7eL3bfSe3mU+sIpdFcIcyI274Ce0BD8ULH/XTRAVx5Kb8kqiF+aurQfKJA
XsR/UbhvgZoMm/1WTsxQvsBUSdDd2KtGG7pEhk0YgndyE7K5iV86KqaGjsQt/9goRLxxHUyiWH99
8eYQg65Bu2VD99OhwE/lpoSQLJC7TxNqYDTuGcH2fjSoszQHVd+0zTXfHWu1Zq0H4s9jPJpjsBX4
srymGk8RS2FrlnJVOWNR6y8KIQOHLXPr6yNt1g89czJ02uS8CorlVyh6r8xOZLEYmg9hyEcO8n+y
KvVXNFwamz4FFhyhbvsiFH8QnPY2XM8jTZFLjJ6wysVyXPY0Bfi3w5ZY/WeqTWkxtB+WdTMYsvrt
Iu4HsIqfAiky1S8BA8gO77s842Dn7D38nemtbHyFKC9xDmsZ6CEP8H+DitXjCHfWCORYP4ReYn09
QMEPA2qcAIxY8fFc2dPmhCAGrLb5M9j29Kp91hbYbqarUb1ejIHuaS7zTcfDMOhlkqtpq0K7kN6a
1UX+avfOl5qwQ89/pJAyRoVKjGieVFTeuAjkKNfhh2faFLFT0SEy03vtXuLkF0alZtbZZMo+47Ir
FZQjRO3R14MkJezSB6IG3TKHHEK9s7BFKUB29Ve4t88Ke45M2dyonQE270de0CrY1DvJ9CAZ7UaJ
fmkt1RnoryFOtEYIZ/faI0//uXdL7/Hz1dCSO3ceWcaeD15rGtDWEAiZAAWvqr/jdO51Z28bBS0a
3BKusp/iMPvfUff3IXyFV1b8+VkKhG0Yx3g9S7MHBdO4W9PK1qMvohRWu3aABO+nZAVS5oVMOqlW
iO7n7Hafe0Q9M1e4294Kq13+2iy2pgZ2HgBzgvLvCV9Q+Lu5GFZD4kxN7NppkEBObt5mlsBFs6t5
WTNj+o0OTL0i2iw5OCOwe/xDQv+SkPMP0u1kXJ5GqcpRO0hAscqol+QZSHRabEHuXqNBKJEzVvr7
b6qSo/lCH1oPvJ4SWn9smNr8l7RpSZW6USd+GuI1Ckdqadpo76oO3NDLX0yvStn/smWxHEx3gneT
w2/uaZy/rBFsrOfxhy0b8seB54GzgaopIQiveotSsYIwQq3r1KBH73tVTwPz7AXMfFqTWgsoLKhC
BX8hFye4vHnUOtYZ6cwbMwVasIxC5FHoXEwqhv0hPcrN+dwcry7MvXuCLGA7ozIBZE56WKPjXdSF
hJmniX3fUClH31iIB85Nvq9UANP2y43bcZAhanrzjgpuXyKKybIT4PVD0fmlULcEIdMdCKQ5WR0c
wM+ks/yhZv+NcWKjt40b0QbXvgAKGkiwsAH9R5tSGkp8H93iHaQ/0yalbcyWrvD1Y9tfDkX435cu
RhY3quCvrmD400hiwxmvjp2DQFYT5+qTIq3KT01DRiKsvgdtFcZ+UazlengUYmjPem7DRpp81+tN
umIH4McoKVRZ9xCMJhuHds3MdjUgxtC9mhojtiMU1ho64SXMHYACc2KGrNG448RDR8LVmIzAN67y
MoZoR0qXw88Hl/ppiifFDaD173AciF4attz4IlK9DIqprn4RrunyrbZ4DIN7pUcWV+lLGj4Y9N7r
PLV/JaD3d5coLPXSbxLaw7V86PBjlN/4p5MG4Fi+fLwJq0n/pMxSfxKQO88/x9jqGpjHpCYGVZ+H
KiQrVgtWGRHb/kgALxG37UmVR3nI4+mpSRAprsVV7XoXmQi+l+QWo70d6C6fYfiDhOQaf4Luekfu
C12Sg0ZuEblqox/O6py1ZBwOJ1jx8fUApBrxcMnNsHVPaPzNCiaE2+3tyO8Ch2WD6sCJ8jTRkbSK
95dhy5xFu9B5wU+TuELhj7gILTXaxeyjqs/8Pi+0bmKhDEgTEYKP2W1T4Ru3u8GGHWt0DfWStNON
et5oS+wmdEEawPg1kOP4pYyDxGz9jQuv4gR25Py2BwkxbeKuDdB0pidtaQBpwFYnMDGFjX21luzD
W8t0MCUF2ZrcV3dk/TQGxnRUovb/PCsouA3pBHa70G4pXjEuaz/3E9LIvQgd6qrfBlGkU9YrMkt1
TeiWzjj7Ea2IFhFFLGE7NKS2QlKprXa68YhD8FKMFHngAfWDfp23+uUhFpI6nLDyrTMfMghElyJU
sMT/8W3ILi3nn2DhOkxTiSa9EXCPLy/KuvmXdR1fctbtx/1YadcisGu8lgM7YV6ss6Pl46PTj6mr
+h3rQe7Lt4SJ5Ie1f6XKmOV/QCtW3GKqpOBS1QCosIm/XYkg3aSMeWf0dRfQ5u1zk3j1wAOtzDcl
FcK33ETheDcoNLf39XCe2WM9ueVNfkYUrZpEX2ULwUFhwKl631fMNryJOT9RmTUGiSRhVptVOBKv
8NPghPqgGLoy6IUsh5lRr+8t68x+KXgeBVMTteNk2GaZfLepfHzgz2VhSy2nHJSYsPQXiVdOE2II
z4P7ZEP4lYrexMzFHVZ3DknOrMnS5LfToA00+k+qeuauoP6RgMyt37VDWBmA7VldJeZBc0sYzHUk
vmoCW1dWuYMZ6y1f7WBMMOb7pq0PCEu6A5pA3w53Ni65mRvuTB00ZiSsas4CRwBG5yy2cod8P7vl
x0jBK4ggm5XXaSOq+NgP/bKZGPKUBYk3hxx8GN9Hh2oax2i/NqfMebT0bGOe5kCHdSO68lRxIdCm
3zZ3ECBdjHqzdTU7ylmoPAzXoPt1h42V3qXGniXkIJeuHR9uzICjRPSOpbsP+nhNtZ8XTOB+bF0b
948ZxpgnNUJvRFrgMb2CJ68ry/d4+5IcMm2BQXVgWmu/StTKqr89VZGUZXSqOJYGmX8t2fB+0TY5
FoRSo48BmlCpgdOv/CkXxoP/Cz6QY105pFKPR1ObVNZcv5OlIjyMswjhotddkwG5N4PqjRNuNVkQ
2yrKFF2JRBR0ZHM00ma+kc5pY/Jhqv2EVCtB1VeytyqRf4NPNlGx4RDe0ays5C2hBxu2WoAXqdJV
RegmMBJ7vo60+D7wbEtQbufJjc5IJ9bTsCVGDXQx391Lmw/Z2KyGIbMwUO9vgDQ/+2bsM/T/2pd6
bfXZYlux07wBgvY8fGc/w3RZhbbvCMClKevZODir2tO5N0edg8FNheHxwfXFLKmS+aQlFRKlvFag
m0KVcFjccGDll6BT4gggpEkOOeBtf8oDP005bgjMy8piX/2r3JvFulF9h/f0W4jPahz6D1fgrl+7
8IZUm8dfF7WVbbJt64pmGYOkKkli7u/Tr9vZvGeP9hvOLDlRfbXxUbuEDrkhjhj8Nhuz5r+jKGSf
zZMZmcfrC/jRr9aOmkfo/s0BfxCbR0lWwlrjox28KjtcdhnjlSwIE/EagjH9TbWo5tONTe6PPvn1
vZRfIekxCasUK4AEYqUwcLDXQbB4L/ry3Bji4I4WbGP96lQU0SvmRQvs14zCXRYYxlHXBxWYw+6G
BRd+73VKBmOwkDC5qzPXKCn9N4rrfdmwp9G0HQ6RYpqtz4gFVrvuFZsE9WO/HEXOh4uFFJuEh8bY
lJrEalEyKLzL+SfXSghuT8k/A5yE4OqH3gCFRA/8ExyVv8p6uZe2SHpm04JAbhpltWfitMrrMnwQ
3RB4c7IuhNtWRwQsG+JpZjq6almra1GK/uzuXNiSGkckxqiDV9VaRbgQY7Sobcs1WLxU2WvEhLLA
ytjRJ1QCog+JHUIVIFjzWlx2YCbb+YmN4QzOmkpjNo6boSIK/mwoa7o48Dk7IEtL6h7HA1BSRi+r
Oh+GWcpEk4u+5GDPm+QtkI3kkp1t7/XKwRT9emo02zqBdNELBADa75vuDJqxdJP0Q8Wdf8FXqTh5
7DD08TSI4emBIwX0TK5xtKuxZQJW2vDrcRD8+hEIj3l5Fkq7/FPjFQsD+RQyCIR0pqM30CXsy8Va
oe130y84DRxCS04FMN/VrKSmo2g2RBe4qcSvQtOUP/1c+Iu0Fas87MNuMpLEFyd96W8A/Va+fpr/
5096/UeuatPcsl6tE7iOrBVZeD/pZVJQw8rKCHhRuvby5vmBAohNHs41NDYsdiVBrWum11fCudmL
LaqJcmuyM/Pjd7TtPBU04RMzv9I3oFIX6HMAQLRo6kaUJGDhJ/65sozuFaldcUEd3RbbjPA391tf
2bV+UW4bq1q6vitkxba242CIqo9jKKaI06cyiwecWaytJaLLq3bhcjszaMGxhR12oxoBQk7LaoLR
bHu2ko3eFFWZzges9axhGGvJmw4GdY6mrNbFMUypjpYR+z/rwUOJB8tZSUyxsCHvV6mUiLzNDwI2
JU1XkCJ0bMx9K+0OQ0EplDSsp0qybBVqJKdYUeiDXZ8A5J9GaWWbWb/JImGXfGAyU/wpzVEJpJmL
eEVNkmRODvoUeB/pn3Tawsdj34S9Mt6W8W8TgSfys34/L37jl7pyfQUv/UDp6mkK9YFSN4XVwGPJ
BSDE4Djmye83aXmJJci+XfS+JHQL1Tqx1KI2BlcI78jg0WNstrKVLtAZQULANUPaSVd1QIUPzErj
7kt43UfHvfiTFvj0P7jCwfR94cFUlPa1XQuuW0WmI0UQiC3/ywjurKU3mofPRVLEmvxzSH9q0tcc
y5bt571i52M5mOdG86mVWk6ZZecLPMFkZceXD5V7wAcoIESJRicBwn72/R0iPzrNmiHlC2wAbuZ+
PFEO0cL86de4Mpiurg5pvtGKFR+BoyFoi38V4Zhv11LMVigHw4Lj4BIJ/lx/ESn43343WvUU0cFn
IczeJQhQgW885l/Z/inkROg6kN+aLiWCh9qVjrbyUqfTZNO2zMn8N3wQKHRMxidEBAjnnppOZ+rj
XeOp9VI5pxrPAtjMBNgLPBJqlxWr6wasNA7R1C9Mkhz7XB2pXJZaJ1GK+orQurq7ZMyVI3S6bk8U
AuswIPPipxYwhZHbTdOTxieMDDDo/t22v1Nkmkmh+p6fmAoM8T2hT+f6neF7LKMfaDM4ypJQ2Ikv
a4OKykm+EKNhQKyaSOq6788PhmVdD/q/LLrnexzahLUL58dbcf8Oc/PlWogcpiNLVQCUcfPMXpzd
R6GJlHmov4BaPNfs4PVmv3a1XykjCEHvlTFFwaeF0PZTrwqYDWQrG157dj4qPflgUqhndjDLXmtQ
vzoOWdmMSM3NR+6GdyOr3q2/0/QV0qXEkh3x9j+7RHBnWj9JNFEohCFk9viOeF4ig9sUPAfZcItX
5rq8hl1h18SwUCLjpzUHIP9asAp0Ht0wTeMeyTbjxamtj+wyQjlgs6hvMdFuplfHskvzzNo63Oqw
paHyk7Y8pjCldSLtEpBd0HDs5IABqJZKNF/OSr5/jAk0/YIuz9BtevdFt3pf3xEj3E9q+gfdop/h
8ejVCT4JKPpBLFfVPewr+FlR9cQ87izDcgtz7ykYiPAgmQ0YJIB7r+hdJkiWRgsiENhUS8sfM9i3
bnNYI7uL5rwUCzldcuFBsOABl2JUvh9dkvv2IosNWRFRUIWozGbpmhPPydH3GHqXh+mK3DrQt4DR
0FEuvulR5UGsJX6PyPGU0Lygl4EkG9eDI+XfKjx3ZiPBlPZcxkIrUEwDY7oDtlcBZl8AM0JJF2Z0
/ltm5fVXY9uj4p/UvBcCE73iDPOpUpOWpTVhpEsen5fDti6t3SNMYxhhbsEAra9JeZm7XSi/HY+6
hCoU0ovektC/LunLXFxuPTpG+gHNwFpDEmOm+q73goZtBx0wYDx36yLGXGGo9OkrTOmc9VNo95NO
M61nnQFS0YOm7iDcPPDQlKLI5Hq1H5gNPWgBxJ1kJLhsYj/g4ATGFuZLL+gDCLiwpmAJqv0aiktA
+1R3mQxlT33+diAxji22TggwheuWZempxyNNK8pnrPCN3bAglA+HUJlaWWyFfm26VQU+QTsIPiHR
jPechn5QZqftR8UVLLB0Ks4fOhlE172hxrhnmYNvAkZdfsI64S7x4bgb6rsyyZb1gMfenQKsiNiZ
H4CEMGFVR7SOu5vmMg0PfSuGFILEi9AhNEZYYapCEBz2nRSUnA/1bX1E5MlvHbScLEkjZCi/ZX+H
eWO9EZuOWDQkCB6GZ/i89JIvZrYnTaLJqWEN4H73/B7MNaMrkSgOByWMRtV7wEMqPOZl1gGZMYBv
ZyTZbNB5vYvvErP2W0jzGQLVbrW+FZaudow1O6lYqZZWGV2Z84QIU/BLV7xfqigpjZmj9touMNEN
wVEbCEqxcxkEf2he0vasBX4kxjJGrByDTI5ilM6r+Q0gn1J3u+SRuC/34Y4nkxUf2kKui089Nu9v
sTkynrP2AWwwU47BL0Hl+FEWqHFMn7iyoi83aev7rpppCeiHks4Mc0LpxF0KNnvu6xz0qvJlf00r
ZSCVMK+6yhk70jUr/AEU16F21C41z8J3p4cYxgSe2nvB1Tc1PgSw9PDUhBfZNKw6cg0MpyZZlomU
HEt1qAvMttI3B+xTYN3mJVPp8vJT0zGtmIN8AuAU5G25JiQi5qIL3SeDGW6S/e1vGumbMehVrf5x
e3x3l73sBF8Y0BrO4b3C1GC+azsfLw+kDyVdEpzR6+spm4N/8ZVYnD5Rvt/gblwj3jtZkvJoGaFV
5cZGkk+a1HBFCqIlTmVucFSycrE306s9e8YspHpe1zNMvf5wtTMxGasi57qnbklYfeT165UWXW05
OdT6q1Tbktn+HQ4ipsp7xN204/DzSGk66LBH3ezG4eX5t4nvISHi96ZLSvL/80DMJLmAlEHE7/Pr
cbzfoOoUfJEzBf2+eIojZFozMDNXmWy+UJLdhUf3TArCR0jjZ99DEiKA+Ekbkd19c6lScr13Mhe3
zw8IKaGbIJuImF1m1GumD7mii2AwDrwsq16QGQcODEBtKNmfzbIFcvtMKMDMM6neMMs7aNeAyJ44
KdoeytB6gXjl2vmZ9UYWf4exAczlfSVge2TVGDsZJcDDrhiZ30aSGvj0l1z3Xs1YnVvzwSwkb3eO
wHVKfOi32gJXEIZmTtddddh54yMvyC4O0AAW1hZ0ReIDr30y5n0Ddx4Pd95rcXmcKBKd2dqpgXcp
YvtXfTQYCd11XUQS3bKc24+5CG0CWCrAdgK46MspzIFaVwVoduU6cINeXnXOxeY/bXFAZenF+j0F
KwLr+ZEnXljfvdhMoSUKc84j17Ea/479SqTkvO5ZEl/Fc5oFVyX98Y+qGxdTENwj97pgUgdCxKky
UWOlpfTm+4pZahdXooJqNy63qSATlGEYZECi0x6aW1QbC+AY801hv4cT7F8+quJdSOjJSL9eRnA3
9e3bbd2/OJX263IRAgnnpRcMIiwuLXuZS04vgR5hPGjU746o4bwGDe9Rjy43QByfMcHBnRE+8fVt
bqWoXtIYEPceIp0829PrEc9B41DPQ9g69HfrxurVjtMMpuEL1eOn+b1XP3OkLuyxt4Qct7B7dC1p
l9BhBcjZfBOsBXpoEg1SrUGHoPplp//PjuULehzU6x57rHk9j+6uoI/BI47iQVLOC+gM51/2rndh
eFLhiFyPxvHCQA/iyBl9z5viWMQ5oRE0dY6IV8zzNe9oz+E12wRsn7Tb0HT++Ve06Y7sK0PoGEib
MjHe7emfC59ZdjqI5lSlb3obIue26xIEG3BMxgzMYV5WNKGdoIE9vy9t3U2ea+gXIelx0lEHc1TJ
cu56ivSMmAjyVy/BATdas71Hby//Vmp9QMkQcAG+V1LCI+Av9sBKGP/ujdGNiVFHFJa5cmdORZDn
6jaCIaJC88eSfRcloSjOYc+0NnAaqS9xz45fRoY43pjHPKYyfMmvtS3niieVHXJjLXVWNwdL+FVw
t9yFetD2Z3/OoHNtUlWkIQhGPb+VeJ8x9UpVwfz6gIUDJ5s7pvXICX3H8pJEucDiP3fnqHEoZrRD
KWnlhZV3J/wbe1UDJMhNNqQt816AGFX2JeIeAeqZfDxw/rJxE1RET9nGQj6wBfUOL7RVuIH7nDcL
f3JpXRsrHGP+b/klAraCd0mUc5n1vtlJsjcNi0mut2nSnZZkuhIUG29WntmeOpi7sYOUv8V+u1xH
T0DxEQoRHMXXq/SY7QKdnjKDDFsXn0ilBFdGpfjlUE7Gs6f0juFHU9hRyQpKI0Vy/JLi4b5PBFoE
ifyov6ZRjYXWAAdUXwlChmoCnXhBJUYQAgtrurIGfq7L+qvfkkBEVCZBF0d+JsJKQLIZO9nb1pD8
VIJZPGfoAtjQX8cx7LP+CT0omJQT8KGHchMSfkOAHIbAl8lkpCnjioLT0B62WtZAUG/Pc7IxIUg4
iwaC6zmmwdALOFmGsBtC69yGaNpKzAu0H+be294+RP1uG6Z0QVo2qANfSM0UZYPvvjwSNZ28cK9f
yPefIco9B8s48s62vdpUIYohkDXRnScAGdJLzRWfdlBdfrlhuvq+M9raY1Qeic8Slem9USaH6spG
eJ7glQFlR189fNUWFXEIwKeyUxh9/ZOPtgKI87L0gapPS2mu8/027297iLjWzqXWGAlhQpiLxDu8
JZJSJmKxxZcyvkasWMMHxORQ23ewRkTEkEggZQyOGX6RnzBTygS7wXv2QEgq8UryNlNvOq5O4fPB
uKjSn07xXzR2aggwSdURF78KWxG7KJKkj6+16H16OSG9dVRmtycRQ2On5viufbBof7wZnHaM2Ayg
M3CMbYoWCQ0+T1qkgyOuG354Utvl/6edVkAr4d8FAjzJ+dX24l4BmDFMET8NiPYe/GSpfhXsC2g3
q5OOyS98i5ke1RCddwI9xZs69mNjIAjqShAHGodRySMuIhw7xerC45GYZ084xPLxbV42TEiAOMW+
LY6Z1zQJb9ymAP9L0EKGoKwG+Scu47dxvHTsj/Ukzqy5eKJFWoA92HYnl8hNfKGGlHUqsRVb8FqU
PxTL6Jm+ZZZDBWdBtSXSaW/UdL2HC+OVjnlxsk1uPnEJwVpaKal3xNwyxM4zLqZCCYWbQx6FiWxN
lSxpyqliqECk/Dh7JS5wkJzgi0LcqU2PR9EmolLYZiHT55ORKyw6aFtQq4V/jgzVTY9tPokQVQwt
qMzZ0cz6fOw9bGd+y2ICLp+/cy4fhk2KcGlGE9qa6IWqjk9dBq8a525apDG2jpnoMep+j1jqjFaJ
eDB/E8q7oPP8tnNWuB5ztvkG3QFDAgu4u+v8vnsjvq74zl3rI5LTVg7a56lHDeDzsIebk8kVatkH
8HY3tbt3MYN9oLVXAA1/kw4Mp7U0rNYo1YjFXmSVyal69BWZDSVJJIi+UddN90HmPalyWnBYoVce
b1fCoyqMC5IyN5M7oDoOGRHDqybJbM610C/VBcLqWgShp2MCaXMWM03P6as0jSNWcQFH7qKTEiu9
DUu/7hfLb8ciQNqiBETdntZJNTwU7HdqeLI0OoA1AJ2x5EPSyVTf38IaRLxcv2q6YyT5ry7xccqd
hJY6y3aAKSuFsHgJcyERNdNZp0GpU22rmb0bcRkjP7Bh8pMjMVZwLP4pLfT+qlN1P+D1lDXRm02f
Fi1cSAjCtc99myqeATKvbwCiAXu/j24ezLIurPEVfj0+GkDL7bFnTLT9mvDfJGVm9gNfaZ4hiZV4
dQ+ZRHXynu5QBnql+HhI38xjY8RJJoMKpphejzuLGmNgItmYvVTEdyOucc9HLalGAdd0RbgmyVmy
/HAHsjJvqWgH0UecgIqVKw5zgAIJpSCUy+9e3yp9gGli+7MbZbmj+GkoXdxb9nQ2J3n/4zsfWCkT
PDAw1yJA1TfrZ4BKCeWimhS51HfNq4YmQlFoYMW/Ojy5ihqUxla6grn0HeJVVFJKXqnni+hNmcon
DmNkKheYnU/St/SZwNAAmuKLhNUuS4sff3PEkM56Er0lqsEQzBxHoFUmpoR2E+f5QduTTAdMW3iv
/QQ6rGeh8p68Siym7/dZQMcEYDgW+N+c6DKgi0GFOLvboRtL+3g9T88bQ+E2ePiy4ExOeUiAE8Vn
5vJi/l3wEY8Aa42PO4AaI7m5nPvNop0f46sP5M8DOffLt45D3uIlTOf6TYXrsP3L/Z1XunjHg34O
tA+XNnzhWzcQA6n8DBjZzAezJ0Ohj6RFfyIy/2szDfnQGfYumVdmdGko9LGo3612fZGVoigxN+Xw
dBWfPgDMbs78QZkEQG1FT85xzBeVDrWDpGwJLIpLUyoR5Rfguyl32d/76Ka/0WXMOscpfXnNmhjv
cKu5XE2+gpIQf4uWXL5Vj3STCn/rhyZcHLAQkRSb6MEaWbQeTc2zn0xp58jupKSOnRc+mCTB5N7p
BUGB1tG9awIN3CW4kndMpvoLYkB1fqcHtFRQHIx0fa2HToSxfMQdtatKhnBdaChrRp0XCWH+n/mL
8sIYMejsuNWkmQBNFRhFAF2LX+WkhNw1g+TppadPdi9BStHCGri4Ai1CHdTBEScm/BRvU03o7mUL
/7i8SrWs6pjc2Cm4FINfNa/hiuS1lu40gCOoPC9lS3KgfVcLG0hFKbsgUWXNo+HrECZvN6k6kTjA
Qtqxf7MSs6o98UIwg/pGK7B0jIjy/w+gT56XKMKzwB96sGFVSeqlsbMtMzXsH/N9zRaTne580ENy
WSONMX6ZpkTBvl7JF+FwUzcVSfjfIzWpw/Fctgwil+VHiF859ZW4/Cl6bJ0inujdJa9+6FoQwNg9
Tl87zF7qMRtmfTmu60LDge49PGQUM/jVU4ASh0sWHBo0eV5kHDuQ+qa2hJmL1WBmSYJydMNT42oN
hishOKrH6CRa0FvYFEYjO0OxlX0JpN3jwqBISLmpoGglP8XwAydcjQerEQ6oJqiyJsbqzl2I6b0r
7YVjtgwK49TnZf8TTkCPmZIOkQPVmmFir441ujGKu56DWo1QZ6Xt/H4aRB/XBF09YIjwSHg3YCIv
8YgJi4AvxdJYdThTUnsxrUn4yY0fmpucgyUbprGb9ZbO8F/djhfpeTZ3ggxyBeqV7jYpsQms9THU
vso+nMDVmQPJnyl/lGtwcRyf3KLnJs9SwZWJ/7FAmzuvVzK7ZF+xLQkkUZOY/wraElO8LJ9RU2EC
DVl0u1+SllHuOMHK105Ejiixu2npTYZuV+olUG6x9J4iT+0oCHcjZj7mdWEu4aGMoQ/zXJ5oiCaT
A2ujtdY/Yijyp2tqm0tLl0mwUPAclOzZLX2r4XPM0eSWYIZgiIhRKsPUMuqgaA1UOKldplJqSbqi
Ubu9CAyZmH6YcNQMLA8vXfZFAdRADo1T3+/8zfi4awArGAYeWhtDewXZ0veC9tM8OYHeWY8Bpwsv
GSrqwAWsZUhErS6UGPCvdghEqoHEZi7repdLGJ+w/SZfg5detlwR6VpUPgFpQ1lkS4CPYJGIpY3V
SPKOOMCQW4Rww3tir5OBXLMzAvqw6CpJUembWdErarBf8pn78coIOBmCqbsSaR+3Zdz4BoK/4uTT
/5e43rwQVwNNTicEoSisqd/MdFnpat3P4yXevgGiI5LkSyEhThNDbiK0A0qj6AdxC0LM44I21CgG
lZLf3LwGjZw5mslQJFm3btfJGo7Ot4xBo7rY2IDwP8k6qHHjwDYRrcDY/JM9HVjk1Yy1fGJUwVOZ
PigqvBst6bBSBgiqvpWwWwt/2csPfSeiP6f+bsPPGWXh/T+vi64YPQiTlUn0u2qx6avsDcaroW2s
EmjzhppfyhOuQO4NwQDIXrXKLuZDq+5nbN8wLli/nrC4SFPu56NudEbmykS/YInFDqSuMie3GHKu
PbJTZwL5ERv0aTEZ+M6FlxvafhMn/MwqYVhjkXNf0YV5Cai9Rpq65hUie6LNfDZ2LuU2imSX/+zC
O3ISF0e03WiKSf9UErcOU7eQhEYFCBlZAKLYxuj5yhUwWEVBv1EOw3pMcZ5255Wt1ZuUzgNCRfVc
LvqiicsNq82zdguPAcq0N7Nrctus22s0vj2eFFi/brXKJv4xfertpU/8UrhBiplEBw9jL+ra8zWX
fJKdqsLiOYPnHFp85orG67g1kW7GatQrsHesawPSodKHR9vaaBT0BHSn+8RVXWA5rgorbiuuJOB1
ZIoQzYnuKSs96XgnYQ3Xux5WP5EQvrVxbpX7y6ouLOB8xgoTCVr+P6Pt9svDI7tNIuOYc+JJN1GH
KA+641O3zM04CqYGWW6fJPJRqytZ9etSC7hdih9HziSL4lA9yY3g8qUR3gFTqNyI1cIlv0xNm04V
1+fRWdRrhXYLni075SHMMqwQkffMhW3WyzjzNxfos+hZolgCIBB3rOff4D0F+TbemCFM2iH4spZA
mmC9PGAzAWOhMYFiuUWQVtluoGoxJISqUwbTiMnI3IPX5uX6ZqIeA31w0QND1q921WJJxaS8o5q3
Ddr5KiyZLJn+2gl4NcECwH4swJIhRtI5VvEN1oAoqV92vUAGnNFc+dqpgaHUKXswJuFQjv9WEP65
sQP5hlLYREQiUVVJvo4yKNPXGx7CAJAFg738YrP4uicZuzJDgdDYvUAuuN3Dwjh+sx3YHSzI5eQW
zMozaxfLFZmnAfaVn1aLxnE3tMEvOtkaZuNQA24Wi8Uht64onmYfh72q7P/xH2EPdcA3khj3tUak
MJ+WIYgjxFg+uCpLK1H7e6k+v8OFZPHBAYx7MfXJNaafQPtlyvtWYw5RI8qz2z5lEdxRizNoxGO4
IzHXmA3o+1hFhsyHynphaHNy76kuyBcihw3uFOZVimIFgvlvf7CJdW2/F1MOMfF9IsFcSeZ54One
rbsUeCw3ZKPS2EwpZhT1WOkrF2RBctB2ZoDWE+N5XKf6Qoh5tXtDYGsM93gUc1LEvIU5Q+SZIypM
F8VK2/a4gJClyVfbU1cTQAsfmwLn24R//LfbR0ULy62rzPnUYhx5j8aMG/kUmmVNgS3gEtsi9f52
7YzwzbkzN9eil8Ja+E/bT0Dhw67Gc1aVacRhTf3N6XRC2g9Anis1NLRdBxbK9tup6Ux/6dd3aKR2
uu4ceNtW/3snYj7XXD/RjZHLTCk0IN1GePIJmv3u5EZ2cCcuGlF92YKzdm9XmZiVgMN0qcpTYhr7
/783IOUEm014VoMs/Xfwn0KdpgWwzdlOKx3XJ/oKrGfdHXEYE7gdWyzn3M232IxBh35GE8ml3kqr
kOzTMRXL/xyEiwJPqUTxUnsfiVElFpnVtRhz55nZVmcTxyEnCIbUb/y3hI8buRbRRF+Z21uwKENG
X6JFJoEX3WzAFBvJJYKxw1CYQRN3pAJOJotRN0WxOyyoBQ3n+ADf0DsshH3rhLw0hd0QHzhaVzZH
7JPUFUKPgyHeDKUgrq/N2t5anjnj7HyF8vHROGQXal1dlu0zbvlBQeYnNJgYH4zoXj65dNmNCtnt
BkYAG8wCyF3W/NXLhjnM8Fm0vsgZcdnABsEh0oDJKtziz1NEqW6W97yaMRzx25LDshp+iVTlsSXz
NQNdelW8bNiJZchdBIyfkWQENjU3QFagmRZ/HrGHle9x1xUGnE9rYve6UNsdSMS7pJLWzn7lhxfh
UlugADB1XLwUYoKm98dU000tQXyQPSd+fNwfH7YhT8k5/apKWPXg8XQjNL7V5OC13V0ZjTN4IN0V
2C8bO995FoziEThhGjH3yU43qj8Yr46toxYknJ/L3stMXcSv7XHWyzoXFLfo0KGCkX83aDsT/ive
+sI43q2fBAx8eapmU2z4mw5wtP+f2hVxdkmi9Mn5NotOIbzICaBKb0J2k2AdQhu2HZr9LVKWFbSQ
GZhsGbcN9gZQKADsH6k1c3piKjlVm9Dch1ofzqAPE297lUuGRwd8Ga3lOVLLLnJo+kW6tIRB6r7P
Qdfb7CSHSLedvyMsTS8i2dhE7kvRAG0YYGnwAV9/Y36vzWAPNbMD+vrRElh8UgaBbB1kralpESOI
XSpXQS4LyKgyiP/D6iJY1xILyvEXHU5v7dG01W3n8CzzAypgc6+TeKCPLZ6Dy68S0Kde/1SavGAP
hJXAx5ClXKYl2JUavSSYAAZuJXDrKZzdwD+kxUdvUJ5twahW0yCoocqe1EV+kx8pcjd9THnLQ4r+
Z+ut2hV54yCrIAvoCnVwwTaynZDfVBrQbnOXFTJgDnkjguQVeRcsrEBP2eMACBOBr+fK+rtjuGcl
kRRDgOvp5poaD6GZYSGooY7HorSiAXCi2iIB38sWw0HAUnmyR/2DsIYoF42ksG9WYpUifOuiSNhS
2lnKSz5jFzELRi96EqmcRaErqzDbjA5Inzc5Ug7504BBxnvexXq1Sf5jU9BHuni+r3WGcrqu0NfB
d7SX3sAST1cbzqcg0iC7pxdoahYBhRtgOrNQ2jQMTVw3vNSTXxQcEO3rGmUaeGnw1I2q3WRormaY
SbJ5Pf6q2jqgMT5NhiSy5itWnp3tA3oqIxFJB6IkNbKLXH3FptgFgjsZChzw9Y7BQOU+uo5AuDUa
LRkZG5lFwZo24Z6oTYznIUODFX0+TjaqVvilE36X6tT+yixnOcNFGu/m2LjN/hjtr2lLyEnzUye1
FT/rUzixMRAhzVI1s3PoJUHOuczCw2aYzAK7lGksJESsVJoe0RTF4NfrlouARjDQIFC4FMfID2Vm
tEaKDZ+1hHO2/hxM8k3o6wvADNk4rdBXUeBzZupEXGwk1zcxWoNJDJzrJ8gMlAd3DLDUq3G62Gue
zMlF4+rPh1SphVOvgAEo7PFxZsYfORqRs14w1xGVt0sd6HLfNDZ1TAEnIMS6GcgGWP5cScBN+Vyk
8j8rdm+wyENxZ83vr8tPuUPMZ7u2n/KlaQ/UYiGFz0hjFRV/rvT2/p8vQ5RUUz7Tbc5iL+WLrLPd
yO3LjFWsDxmKsiAmrSBFYnSwtGBADMW04tdHh6y8j4VVO68AFRB5vYRefTMQlcxtMrE8PH7D/JX2
j4Dgo7yMC4OJBSbmXXrEadfI6M6IV3y2B4Qjdwm1hI0nBtiBVHqPHAYYrdPqibZJsfG+j76U8i/Q
LBRA+vhEkAG/lyBtq6C6MeeBqSnpj41RfsgecNPScG2JzVjofmalSZn7rYruOW5LSEnZpwZSeDPz
2sVzeDFDQZtTIhpjhQBzr0Lk8xBTmFzE6uVZGfcEIvh77xlmBAJBCF4+L6dJYjvDdDaA15vRIVBB
1DcPkIRzXl2RnXx5jWQM5jEujA/GDBC60gPZD4EZ+ok50QNM6fpWgfxwJWfkVVnquHRpQP7HC9nl
bB4DH2XN/4Ykb4l3pk0n3G2txK/h+Oh5jwP1qjluf0ftWJkOTYXXh/QR1SWzbzqycaj8fFxIZfQH
0g+rR4t0I8w2sue1I2qyNuhFo4BeSUqQuKOIK2KQURk9rvsAsncb3GhlRUhw1BtzImfg35IA75in
Jblym7FSWqFcq2cSBKV2YbewYbx3fzbc/Hhr0CVSxdSRqjMGWIt764YFHY7FfwIXsz9VKkmF+GvL
s/QMURXM2GCTVmMt0qdkPn5QydUwk4al4BeI8gfvM1f7Sha7sF2XkPqGD9gxRdT9eHwyDNETXVgQ
TSyVNt5SccjhB55f/z4klV4jNCKF8JB/tA00weDIQeLqQiadjsHT8sjWQTTmyGC0LHL5ssf8BkZL
AQvhzkpOz8CH1+aVRuoDMzlX5ogPrpbWmKxF+sX25qpsub4I84bpF5S5tfF8BGp/SFE49+0o6UYG
T06/Wug437SFvQrgSA7jf7DgMrWSvziW7Cc9yFVbsshSXU5VArUAYcId3QR7ApavlpG0oAR+Wyuq
hzCnul/LoL8Ll4FQTGy5SWPOR93ISWGyUT7Ex+ex4J2XuAnbCEgJPTxCj2NoMUMRGoFO7UDgI2fW
H2ACJSPwKGWX2z/gZQSDni6qakLgJhypLm034128YzRnUUzZqvqnFUT1dPWWYaC1omuhRDMuYYzR
L2J6h9tpPlSwtTBh68akFRMk4qYx0hGg4o5NBjQnZphaiHRmAkY3SLiL+bSBGLGiJoi72ZubjekZ
koXd3rHOhNnLl2778D2WBwplpUGyyKniZQOACEGDIWzOlKWec7prX89Hcup5GfWFQx07sXo0kqs8
TgeW+yPm5LfGVfBNhI6LP3Gf8XqqP1RBWpkuMHLI5zC64/uZU1WKHFZh3kA5LgQU7poi0CqA9LU0
ZxWRgbmhXp95k3u0C5p0Ysp9Eb3jWQ6a0qJbR2ogBoU72wgYnwKHexUJX9sYaWnoWV4jTrbQhAMD
20BRLrmFZebEZi1Hg/ImZcKYYCXwVAkRsHIYLM2Qh4VnN8inHdaKk3wcp/0sLRVgPG+0mm1K0qVT
dJXTqeYLLzQRCaLjWfxaXg4XnsBNXLdeX4k3b4ev0yBrM6Iv30WUDUwrJr+FAGO3A0t1YQBvTWnZ
a0PIgzNhI2Cc4iJotG+R79gsF7Uu7Kj4DiDaJfd6FMQaKQK3WHDjKWncmxk848PJN8RJI50iot0y
QIECbhKLyA6Pe4Gy0wGJY2aJNYhz7SFuQUEB0RziAuPLMkD3tw6Tfk4uTMxAwp5ZNd51lLtiZyvl
4FUOR4gSc/mWgOJ3wT6Ue3OoE7G88mnNFpJ0qM+5DV2KnrX/jNEa+l4G4ndK7Trh/5CEUo1p4CzP
IYJjQhe9ZINnICrscrI+6ztB34RvxiOzJCtV4u4iSdRPYel+XbWuqOn2KzGMNjPF05drAfnFnoiB
zNkUz6PHRbmkE9viftZlv2kbxTd0EfcyDil3A1wEPTJb768rIyZ+QD9lyATuUL/hkumqEEjXDC7q
bAMhuXFAoA0oTNANSUt9NaXjLBMDLlfi2a/3GVm3/esF4Sh30qhAQrX3zVCvJvIa6jUQpnUayHE0
6SLxvKXbZ70uGP40t7qhBSJSOxp5LFmNRRXjggr9IHvxyjMy1zpEfhVvz8ZNJ4Ndyz5owuVKcgvN
75FPsNXb3W7dayLRyEEU+Zf7p+pxD16igvCHRtq85dTVn7K0SBE6AvuGsGu/SVNX0hjGiv4RVYac
gFJw9Upgulw4G47cVDcwaDSBBlE+kpQwDxpCnAQJ5UZrrF9ak40PKJfIAB9Y9333Z6JtUb5/aTgo
Y6ivw3mP94UZEdtcNiDlbUHl+LABaexScXINXuPp8IleR+lqUZlupSg9Q70ks84Z7Yqim5/2k5gZ
xl1LfhWWQ1A+cWFcvCj3cM8oCsedzxhw6/s6Snq0GLVTsezWuUet7dCIYGYYcjnbPnu6Fbp3QjXm
HRiYXx/h/uELx+HxdGZjB1/3uKdNB2QsXy7JSFcZKBP4W1NiZQDV2Y9RNSbyqhrde8VyV5rmE6KD
36gdkJkhiPXjCSsqq8Q0jDLJfSGgS6yZAtX/+orBwh6iRNoPz43FCE02GcC6DXChfqI52tkcpLUc
fP6x1/Ni3UZXX/p74JRhjoRuIimj/ak8BkuPaC0DhGRQ1S5deReN6beG+xTAyMjLzVozrAo9GpAV
XO1qENqZKkDRpzYKAKxYnvFA7K94+uFFMOhblEu4SlwO4QOdPfD/I+2BWVaWlROHGjIeptlZR5d8
ZI+3hci2Mw2la6ZIGSmES2B3E++AJLRi0I2x0QxH1kjvYHdp96u8lIqNGhfBC7v0eIWIZt6E2rFr
RvMDD7v550bkdK3KTSvnsNLXcOF+S78typfh3Y49cVJbXDGop/2oAefcAIbDiCOEdaQo4b3ipEZt
yLgYXhIs2pAlDnhu0k8fg1pVRmLvlml3FXrcEc6fvkYqRk3U8kQl/vwa3SP7esAKO+jvpZGWxEm5
yJVZCBdyQ3bmORspUVfgVEESvmylQs/iZyyqkP89CILCZCfRWuDthM87bt0XT2q0YrXFdj3jPrXe
K4s0NKICpYdiSmHoraak8eY5wqN/nRomBWaoggYJXGasXCUBH7HnjOZ8CT0lryObQao9G2W/i2rS
yaBTVMDTSVLhocgZTa87SMs6NApozWWKVIgEBThl8dP3JwIlS5FvyH0oz9JngCc73OmcEJkACgIq
s005CLokwO2lKgjtHSTRpabXFIFv5qojDc+XNImi4hMVtZop8USsZqIFY8/89pg+m6O9z7rdiyri
m/hn+2/ID3CXh89UngTtJjFJixVRPYki3p6U7o763ZrsfFUDyhaVJX7/CBduLet1wtk8Utd3iXBT
WhNEo/A60kUaUIjQ9RhO10MiznAE1D9vk4xgM00S9AOf5ibug7uE31prPuar3C4AvfSrZ2q7hvJV
4ld8xPSsCK8QewzsIhMjRBMv3A1w4Ere/98BeIqcp5Ujfb9r8O55XjluMlIZqn20MUOjFCMZmQnY
gHeax9GYIsyxaLjVTP8sWqdkPQi6SsR1VQ+MZGHeZ5E/ij7NDDQb9D2yK2r8YrOjIUHKwc+CYCOd
Q5ujSEnbEyqal4R/zplF7aFxg571IYjggIjii7bbLe2TyZEdBeoJhaS6pSMuWJlXOvwrahMYkFv8
1DmbaWbVJIN93E+pDQqxff0Ls1OQSn5iY4QhVCbnHTzYR3rN2ptmxijItlcmU+oJcAP8L2m+8VAT
1BPAlwV+aoRoQVNqD4vTbWxaH/edH1jVR0Jc9L6Y2hDEBScMurt5LLTLn0nqs6ILjzO9jPO8Zpjc
BA5msMfD8FsGDDAtwDISRxu27pgoyufm0rRJy8ZL4nPiBd+6+HS/vcmAVTxLZjA0o2idQ80YZBS5
IHq4XzGs3PGKdCR5BZYwg78FwYDU7Cj1IjitFKh5s17lprctpnjRdQvWVKEOo9SOHXTRkOiy006Z
m7+Aeby9azw+KILdhrIEMWJgNPyZjaaQ1xC8jqnN5mJiUzDs1Ng4g741pzeQBCTM7I8jU0aHcd0G
pad8hw65ZMdDNvnCRx4LMbBAPu7NYASWkxxUkHeV4MkvLrzuqeRxQuyW6o/VaHf/hs8p3wTIpSpc
9Ny6959vDwWVRe366JjRnG3rBwv09Q9xxEoCSyEFUTDDKabuz5Vb65z6NJAwNqufWOfN5wKCRPg6
FxnsAzgMskoUUxbaSOBaSw2HdiE1cu3xX3MTkcndrVOJvqr5lzJoMSmQfCw3Tbi+KlYOIMT50mrZ
Ul1oUCTkfclN5zWbnKX81zErwgyicPylXYIuxrq7khmICwU2RljYE02s9FXeI5gNG/ChOsjQUo+6
LgPB9Prjg16KrrPtotw5myFK0F6KT+rIRdoi5ag3XVnko4qXLQr3s86T0jqSU7/mOoJPbVD6LW+9
4poyre5cR9NOViE5Dyj4v1g2V3rCu1gXllMvaS01PLA6COoVfLpWd5EtoCQaFShlLqMuxQpQ3ipg
weeLvvH6L0wjVMLV2mwivvY8BvB/hUd1GdZ3KgOBz3/Kx+kZJMxIc5BGjrqpgBjA5A5hKFZ8PpYv
H5VELrH5B90NRjXAJZeVB07S63dy/LM1HPCEAN3ipWJ0ihDK3ut2mb/6AZxQUHlqm6vFSCADWbhi
UujVQfljieRn6qLnMDZwTOHbV0L9/JbCg4Nfko31mQhE09hpNFVbCqzNERjUQvzagn1Gs0gW5tdg
o39l6p/ZbUCjogYtU36vT8XcbGJ9r8A8KygASnc7aj7HxhNNDlQcrs5mFm7DXb1KvVqpBq/qNbWe
wytiFdnziwIXOlAnwpVyQPW/4R4Eg9sqD4iR9LEHrN+EfABDS6HUCxKW2ZVUYbv+lKEMRUi+pzuJ
jwNS4h5BjjtSNbLx+iTqXQ16qehWnMrQ6//zKnwpvKYqfiMQOc+rRG6RIp/52RTJtvJmRpWZ5/PF
OCS4WhQHthnUnCDEnLJTWCXscwzl3Xo+XetyVQApJf6I0GT9rZU0/ITyL91V1lfWHoD3dT5tldHE
V/2ppVKP3uOZP0atfLfVtTNohUooW6YBLp5gReeYpI6Ibn7v3m1tJBqfaKIpHgFzUB5RFUyr0e1z
772Eupwsy8v6CiMmDqQcIUzuttC0Sz1qDFM7JoUcuTM71eHFAhGIqb4nGnswXuS2Hkzzbu7nk7fI
MuPY7A5TBR/U5b47AA2J71SMPCRx8A+BePE0jCW6WYuZTmiasvzkMnH9GQ0DQZ1g736sDzLOIAgI
DlQAeU9t7opSk7HqV59RpFBh2demYZ/v6l4rk+io45zFuvQWx2YVCpgOnlhSgFhABInlJNnjI5PQ
Q+tDzaXMDe7ZPBLEPZ+OjgLJi6jC80T55lBAJrOtGfMMrWICvCrZZfE1DNGiBDAjEHg/BLG1r9ok
9BmzUpr4DcG+POX/Etat0UcRXdvW2dDykFrwh7/PCO+1Q+XhaMPMHQZ8OVzC/GEoOfdG7iLg77/x
LzVTddGyNzkOMKjtD/j2bOs1vtfzxgNgw7tfWkLgLFlzauPiS8s1THAWqXi9QCRCLp9OTHHTAaLA
ZZQTJCzVc+TC5cN01t+ni4+REhZPqnpXaHrtCmS/AQwvQ1vfvLt3wO6PqTpyp5gNUwMw31LaZ04q
WkuiYNlfPop7iJJslOJX8mmL3GC0wzQdnhP56gWAe1KDUz5PnWxBdBXA5v3eXizAlI9PYittaK26
PgMlEnCZaLAdgeItmEd7UXhDsHq4eUiMHYFa9WPmRXUgH4xYvmjUEtyYXp9dM5Ui2IK6JkTwO6gO
ZpYEncXfG9gxAVe/s3GanFsemS3MQtDxe4ecXgcM/vAya9B+myaY1j5UYiRf5RmLlnk7aMdOCgrf
90OPjhi/7kDRyRzTKTBEQyMaCkTLE6m3TGf7+b7LLxPnR1S+7m20yNy1g5SBSSbAb3AgyqRAI3ZC
ZrUlZn9C8ZR+xGlJILcr0RkdK7AwKwNy5K75pDPv28zFyHhRwESVlnqDe/EKWYgODNs2/S3R3+Y4
/Zp0UPaqJx58+XgDB1xfV0+0XFg4xAEjBvZzA1WFzshX5Yhwq7xVTzOs8OZ+ZFF9+S7ZZffIiDM9
Bw0hO71iLXd37WlpHoPlqmDnFjJkAuX/CB/DRP8JZL1RQRyKzc04vzuHVqte6Dfa+iZnL8tYtIjP
TfIcX2bCXPocCncUyY0ojt87ukkBsk5e/uaVPNIp/sRfVRImH8Eo1rB4EYda7deTv+XkEpfwfU8E
SgQWCv6PbKGksBsVt0C76PzL7Gek2JVMcJz4OYbJ2YGhbDawIitZg/rbvT2RS+cKoTO/C7Ssq0oK
Zt/+rTm/KLNZtZ8eb1EWLD2xiItDRP0k+p52LROWioljVbr9/Oy7U2fGA2HC2XJgaMQ6zkY68r/o
XKVUFy8xzCY6oQU03P04W2FCkf0+LJtPzKp6uJDeTDQWaeUKSyeV2cX9hJI1/s8k2vkwCx4nX6Kd
9PX/q1WtjTPnOBedbfuU5tTy6XrHzRJD+ZTrZEY9k0Gf8BeoKqQLz7MAqP5Ce/WV5SytGvPW5d4B
BGeyakMY63EL9mnR4HxBvnW4xedw4UD1KGh4hAYvf+JQqKQvQ90U5fwtFbdFfAJjjhNFl8l3F4Oz
0ij5Eeh/U1SM8U2O1rTI1ypfhZkB/1gY6Q74dU3mnMxP6pYpPtUlyUne5V4sJ9wXHS2CEZY4hb3a
/kCNmbiZLVHWGWzL4b+eJHdKpkdUCMnYwRGaFzr1/KLdQKzv74fklPzVCrcE/7YeYM15qo7Zstoj
Cc2nftBbg1ih3R5D1aUQopYu50fxnZtEksDteatYziKMGM0vUzY4+7fAYranPPClD6BcmrKD65ex
BxpydnI/xrXwSmq0nCa/78JNNa5vHXmGaoAZqpxcgOJ4cwVw4HTSMDYls2iXPEiCTGXiG5ewhqxC
kryiH2kCBQI0N963YAQgSIZ0wEnCnzGFWtIcorKkooDvJvVDqgPgba8u6m5nojLLfNKiuvSOVhmw
d3nP9npzVhDBN8Mx1L/FAqaQ+a6chOtXDoCtWyj2PAIhZ2JvnJU6XGGLzl1W2o2eD+hfU3yCav0O
C71995QXVCiQKaNO7c7jU7OHmwgxZBiDrpE533oN0oZQmwX6S2QUbboq5QkipcVv1aCdIhU8ebAr
l1greZbaedoYO7LHaIIuTvVUXWRWGWPozq7xEPRO/WaEPCY+RXK1OtPMyl3pysfuwbzby7OA1SnB
WGtWfhVgyLw3XFQGNoAg2MqxT7ePNQxKrba1Z0EtVn9Li1QSU2On2DPmRJLmbujrA/DAavBQKjxO
DnzY2gBu4UICkO9dD5sGpOmqtB4JDgkkQNuN3C5Ft3dAL0Sc5IaHIXXw71RrsfdCB2QpvV5ePMqx
nzFx7p18E476JXcvSTuAX1DHwgA2a+qB1DFVdnwUSvYWWVbHa5z+WIuUyfYp2ByLi/VNTxpxxwta
12LblUTGrirfSRhohsRyWZNRXFmtqzk1WBW/z3Oa5kCGv+yjpIbi8lKXbO786yu4bCpjF8FJhRU+
f5n07zJ3Bjp0Rl8eZo4Wad6CgOLE+n54BG6HWH2VQfpU4aOJgliLdQhPG6P05uNjXrRQ2cFUClfN
Tbw/dwO/MpiFexWYm+WSv1Z94ETxdu5GeI90QNWUx2Ey4vthWV2vgY0jTT897lVpn8EGBh7Ck1/X
dr1JGmYlbqCqs8Mq/VwFZZlHMa980lNyXKg/PaBwp8YKqdXlWeDDqPu0XbP7RPhU4r6xLExNq0dI
3lImay4nMTD8eXPBImE3D7inJMExyHR3XBXrS5bT5F6DvKqafm/lB7Q8RDYH3AaKra5xvULCsWJf
4nOABRe8QOB/4/FrBANvEqI+afBJjsyJ+tSPAV64vOHHr4GmSmZ5DXfKqcTZJfyX9H4CrD40EOOU
VraFPIntoTs3g8igvR/apDXhMsjvKc7nVzfkBqUnE58J6tnLHphexhUo1AL8REI43yzJ0kpHGKu5
ySPUYUS4gq3OKlttAbpA28Gx4hhr49J1dwcT+3xUnR/HjLkiYtGHJS7706Z/ubTClE6Z80RO8WK9
47stc+GYqE6QC4YFfSPqiz/iHQ+m8s6YT8hXLVWFeO+dGgrAZM9c5W7rlpoeOa87D9FgUEdliBP+
g+RGgqqZR4CQtyrSiA4rHsDGIGoer2PB/JwQaYylV6IiU32uZrZ3nb5gfoZWWQvOrhQJKmwRoFDS
GfmLH0OvaMQJC+6g7OpiuHMRJBtUgnwGjb0WVvG+/vvQjoAe52SbkFFq33cMq/FqCe6hCdZlVv9I
F1XNwSP4p80J4VoVT4lVG34dIPpApOy1VD/5ZyV3AYKDn4eQ3A0FyNl9wj/yqCawJ/zRQk418Qqf
h5cHzbhUCoJ/tkCrWzm1Tg/gm21xTsmVUcGcNzZ2PXH5K6GlYXhjrsDfTs8NTVk8NtZ/awOEX1ic
k6r4ArbCtBb1CWnK7t1Kucx/UweS1HQDQDv1wKPO3g/8THUGXRJcodBe1FM2omQlpG7BnmNzxMPW
8254aVRUrtxasDMJisDmXd6WHXycAUPSdyj+WNJvXe0bwlbyDB43IXFnEIF4N4c3UE7RqN/Dfhd3
zadUMa2DqHZhdACOI+95fyEH1pJkEUTYFejEQV8B39yWeAsFP7G7zCmMYG4YP/3FqsE7PQ5lMH6v
lsIyaeuOzfSKmW6VsLhzhJABEuqnJBz0ua87icEVUxKURe1az7mcS3OV1jwsXcdGpdlMpovkq99i
/+Oj0vLEWNyhZdIFcOcSaHAnYQYIPD9EcySNP7RpLWv3be/ONNOugT+CR9WqN8z88rXEIvJSB+ix
fZnho6c5VCNzU1dUD3WKxavGwfERr2/1nKqM7ZiGbfdylIuCv4iqaLF9rLZL1G8ad3fU/bwANijd
p9BerkllZRz2Cc5sz4LrD1veJEzkXY7BArVPo2X/WZOh3NAg3fgY0YfBno/xZk10PR+gA1yPYPZQ
a+0xoiJ933qRw1PeB+wKNiyBABFP+SLv7fl/YoN+z8hC1AwOPvrMileBCa6ujcVfTjeV9A+LZyjz
4d1Ooqj5vg+5ora6qL4m3nh3yr88Op7gdRwmONjatGRQaRNYSQiGKy5Amu7uXaheF1tAfsIPwWRZ
GVBgnR8WpekdITWymC2hBpmT9ZXeixcizPjJQc4xif2YgwAAGpkudf7Sr4vWlDur6PxrpjLwBBrM
Iz4Q0JK4XL7lfE5LRRg5nuHu5jtzA8vpdEeND/Ji4GhVnWOLALNQS4h3QrMK37hB8+xVtIbWJ3kF
/JT6CRzGxbwHMG8P//crhwbyj/iDO+TyrtBigQ+f4/2N2A61zYQK6/r9qnDJh1OZn7NluUBGN9fu
sGTGzQelS3Adrxbe2VFF2t4KEY+84rlR8k5YrXDOPAqiGUlLq3xYqy+Bi5DmwCpa+pYjakSwvJmf
8BZ9b7YxvaZw49Gjca4waaJcUKJwmTaG8rccaCXg6F4AhPkILBKNziE9XMnTBCiyfTSK5K/olQjp
t8ft9Wv05uoB23fEI+U7RHYnBw0yauitUi5dYhubhLMxuF68XY619aVNMbtt6c9dXoeiuMcA1u0X
eUcj+T22jQlKnLaOfLAINjVa6way83FapaGIqhkopVhFWBWJWb5anewIiloCQeF8y2WYzP/31vUP
ccWmq1hd8sD2yp0NU1nZhIt54L4AhO3FHfEfyyLouNp9YChCorQX20e9NH7igmuzAP+Icy/+mnkw
6wL0RyBKmHlHvDhRK7CtXQINcc/lRgPBC7GPhSb14bwPvSzcJFkpwGhCSLAYc/Aie2qUxUurUUE4
NHdxJp0sBFDZq4OIn3SJgWYwpGUMgt06O59ZkkbpdMt6xIEGMAcYrQVr9vrBqUNNHbYDJGdm7BRl
4EOnFdS7nCI0yBnTopROub7yaru0zbXq3TU/Pyy6UFB1diEz54k8otM40zUvSit+g2NMxKRnW0FY
TF9Wf/6AB8GVxa9HEQ8lZCtE2WAPMTkS7Kr1KjPRk/knnTHmL/z9rMP/BTuTqJPuNAPXDRQi+zv/
WbQMwUm4UPMOujTPPiEgdCbQ5fqEyvapLe8O7AXUqoBH+fqhk8paSgkGkJkpVD7vn2dLVphTEduu
1+QeU0ylL4lbv7UHr+pqS1iBGXmG/E5GNZb6s6hGluoHPz+I2jCk6DDtboX8c2rGX1HE64yZuiBn
kYUl9rYB9+LIGf9Rv3Pjpc04dbdQ0QH/zC8xXg9Jz4gxMgWBi+lr71XTXgpTn0j6Xd0xs69ZAoP8
90oR9aZTzqVb0GwxedaixpHvEyjfPtpqBrpgFZgheFGBzHLh8vLZJccKaQfMW9TUxmLOmgU9uxs2
a5qIUZwHfBwQhVaQBnNLMzrwj0Vho93uTnFZIPkojxrxtQhNooC6ZSXs7YKwDpEtaldcKlPPWaxn
xpBeW68tb7mk4CCNe7+U05d6sbpPrmGNvWieRFlNODWzAICyqWSPRRhknl3FVCYfUKcu4he7rWF7
nX8Plk3QFkXg4kYsFY4+7glPuh8YOkegEr6irTNUpABQ+4Iz0q0dulGGI6b1qHaM8GkIFzg3Hx/D
BUZUat0poYWLSpTw64Pyboh5MhvgAKy651D808DLzI3nrsFqfuoROYm6B1/yiBmF9QWNlLBFGXYC
NEmxrC+prKu6CUwpLarMHjgojxqUon7WKLWjcgP7vKJnwZGkcgoqzpy8Ou1tOWhY1+v8SFr4uB9b
043cn+crgnUjVOSQwqgZ4y+wN/oOnbnSEPz0OaHY3ykclNYubgYAEoCXGT/riFGiq3GtTQVnFBP4
c5gM2C8CSoEtj2OBpQLvO8twtacX0fDENB+thq8tYyBzHfWhHJHKfO6woPK4Mx/ATygy4mrey0D2
mlqchyG5wMcf5mBwuFz8sdEjooL0CO+xEhdj86ap5AMhkB99HB73iaKCOY6g8hpNGQ9xyvbJprZ+
mnGbIjt1HhldJr/8P+tQOkpHoxSj9WQqOngQ/NV/pDcAfHdw8Qv14AuPyTi5cIw608ojzpRParV9
LDz4C5zHImic7TgEWNSjGSVvigoJvFAptoUnHh1Lydrxuho5Ss+MWrWwvfKt6dXLpJzkop6xy07i
TB0zuH4ytuamCszTSuzfa3seBThPa5TJrCggffVc+HagI82ZTTMfVrdi+ozZwNetQY2bQh8+IIDL
+cixd0u+1u376kH0eBLap3EgIzPfV+t1Exne5HRGyq/q629O1Y+7+uoCWpuXpqyjBULXnp7SjJ9Y
Sh62Pgnhd792TxCLeoqtFq3x+s8pWny/3LRTqS/RRWPfTuq67/sz/lZqXShgmTrBqVJMX8GpXNdi
tIqGSNU5rPngN0Asbj/NdV2ASWb5LWrdeaRFoP1CL6yfRySOXXnsnUXhPvLL6FESUApj19CxwRj3
5Hepyzq3OrlLQR67TkWmjS82G4ZDbxGC1DefUJVEWHvXwpRYHj/3hWpllMbUYFIBurp8fCa8OaG5
nxFEdDiPhRAobPL2tyIkan4vSTGcv64tIV0ZNNtlQmw9ri5IG2SUyecaCAWuxNPg3doF5hkzhNyP
F4gCrRgiN43qZ2uB+yQO/uLkpjPsW6foanW9BR/qnPRnt2IJftCYExA3uL+gebDRVfVHNBCTjOqq
eNBsW3LW3Q0iwluxxTZfdbgT6m/wHERUCOo3TKtGtQBl61o4BZmG6hUylXHfCs2zoj4oVoR56vEZ
85I4WmvW7YP60CyRsMuq0SHYXVZATvkgJAj9Py7sTob3/S5qp5Xe4m/2lBB0LzyDi8xzlZWpgHdl
Y6EJJhr5mUbdYxHQ9Mb1PJ2q6cueb2wRT6F0+l0Jpf/vR558mO5FtYwSISRMyWHihv1Hlxmc5iYP
pfl9/i++zronzhs6ZaCLMBZ6XRUwDWiXmRcTMGW0LRTxkXjWirOY0Y571d7Xt/cDMMPKuK1bVdgI
p4Occf6uZ8l2vJUdvptxEODnCBpaXQPLLzu1Y4LCJPK6cHAv9yOeW94xDHcXmE+cbivfqH2NJLwG
z7NKjnMU+0z0B3KvGOF9A68xRqOl4Kiri0LMEDitnSJs7cyh4h2BiYrv/Lu1PQH4FTP5xsWNxbmf
kByrJmFsDjbIR6E9Kd0GLHlqtpTQJGy8Sm1KdxJUIABQLaxg1fjkOXcGsX+UNacnyDOg8FLpVd1X
CrJ+uBC9w0MKyBW4tqh7M4NYYhAP3mywrDYqpXxjNJU/MYOJ70Kp8owu2JN24xs4Jgr2t1YCCRFA
IPoR4tBKlqy0dAfAW10BSIRW1Z1X9A4IQiaYvg5vYZVxHmQASkvPwZSWVYLsAYLh8FLFIN5sfer6
8k39qw00HHzlshie3I6sr8Gg5SAMuxBTYiBV+h9qSKhJFOh/hNKGUI4CaPEtwoi0rhI5fLR+7P5H
UAb9uwXI2wd40yldLwpDH3zE8kHygTeMtAvPq0oqa//iJNn3e5QzYFhNz7z7JU2XGIuUfodbjZfJ
0oec8Zb9YBiKIr0cJMUBxJ/AT5KDT/Bzgg3smrM3o72ikzrDsh+tApJca/1wcaG+Z1c2M+tlHQfC
Gii3hobT7qnAMeMPB/eAqHqILYrE4PkP0BArg4RjVSYYN/GA5R8m37/U2Daj/0gWX2eHaNdQS4hr
lQ1/M1NP++li2hu21zoa15uNcGB2GjXXNdMuC6YsJ1pjuy5oknyC1ozQBka6npX6wG8GwqRDEGlj
lCV8NbI6J36lanpNU/A9/1ctlQsUo0u0EqRWK3g8B9UlyVNgO+IHWs0dcEiHLn7gzErxjWVR1K6n
/ffFb9vaJYncBm+uwlgkJomUrVnk2o88DyyLEiI1+Nxu6XPkEgIPj7IVfJF/+vBeX+DD4eBXy7To
aIN9zsSYGIm9qCp23bqBIb8ZiQagfeYj7PsJTUQhpRDeevhmKWOMjnuv3kA9dtRzpFpihq8lPK15
gZexurKLexbxa9qdwzWb/WzmWbxASQecTlOsi5Qd6TpntQ9OUKEXD20VXq4bq18aBrNYElZWSC3i
ZG+1x4jua2HpwcdPpyLgyyqyjrFZKOXe1kjVHcAhZfEhKqMQyka/qPH01sODbRT3lqb/t+L0IKTE
Jy16A83bCxid2hqsuR48nivki2EkbLAHfkXSLyolK6UL9vaUaTno3Vav3oDNrmBypdlecci+2LiV
Rak3SixugfZhmGUtYZT/zFwqklRDoJ1y7KyPUSOC6UmeFHVz8ASFCQopHLM/6P6bp8rGrDY4Kxyz
he9fsogUY8IRs2RnGwsdFTU+YmqeHeg22dzCZGZ9AgaNduNLurxUkVoW1/KXCPVQx8gR+6rWtomm
RhF3i0lbEFWwH0fXIImlWO0MvNO8TgOYNwRrvUG7n5aJIxBgIVc8VvSWWU4DhORTEvUdv/+CNQUG
kahEhwUQkM8N3KX9rM4YIda2q2eOAszAgDgtSfWKZXFIHapiBaayzgT6CpyiZ1otT6Ko7bNFqB/t
yU8/NiDBE5DjGgCVlsRkPIpQYtzJQ76itFqTTWbBoP8SGmROe9Udi41oqbQazRg4mp9a2f94a/z7
N3Z52OkJko1vVtbaTYK+jo/6GPIH92buFAIz+y5BW04eR41D6DZH2Qwciz4VBCJaHUk/mhluhbj4
qQ64rRMyZsBdSWyyKE7m+bFLAbdCWCEJWHly2IJ16Q8bSKrpIoobY3C4eidb/2OLePn/rlwSy0KB
WlblLBEU8O+DImxAzaOONg+AOh0pNOK952wmV8chE5BYRaTMIDSZGRyiHd8oBPjU+eihJxwEglz/
UjoPFQck/qeQNjRfkWIWC6+D8xXR5Yae3oGJb3CbltNomHwYLaXWq5a32WPFbNWGwXjHVSNpmPbw
AlzPUP6iv41dWsnfqDuBNzvr9fztenbJcgcf+V3OHJ2HtmI+1FmzbUsX6yHJfk//i+XbL3FednlM
hhYQYJrDkI4Ms+CqqIzvErErBSb78CStqxepJydmnTsroKSKZAEvAUCea6ZXDEu0gW/0IHHgb62i
AhA2zohI25NPSNDmxfUqVe/eLA2jie0uWfiibvatg69dE79cmDiCacnZ5X8yGErf+fpHikVjTKyC
BFdvsHHmeqoxgLXdgTPL+pgeb85MaeReM3NtRyFSplz4W4Eml6s41CyFqp3IZ3DnItjZunjU/pJR
aK46xjdJVB6CO8Q4Y9//ibdED6UGsKRrX51Isc5LufgVrtzW0aTxFxNiB0H4/5ABh1EYsy4BPFLC
RyLdXzrvXovvd09gSYg8+QrQ82sEoqokSUx3Hg0DkHiUAHcFcN2uM/LOsc1/gnFIbTIdr3QDaUmt
nHg5GVZ8mJc+DDSTFQCypT8xUec7tCBtnF6iEb6Qv59kjxt6ir2VZxtW7hLsilKOkQb8/l7GWNsU
QUwxsmMze6vfdoAwoyCY2b2XQGjPWJsSZY33TLKwo3Haeye4SKByWSfnj61iK3y5cP6Bm6BvVVBv
Ca+/5noV/55AAJKGoBFoKaOGUSwXOPYWgl+ZaEL6x7r/2VCgnwzks5srcQqduEztW85dh93ExHpm
WjUiPZyW56tfRAh2n0EUTBf1UrsZQlMGnd1joZy95gcP3QYq4olsO9fat2aMotADTkLjQqIjtj32
j8D0YDJlpNNhDv2VRGeMYTA27VmIMjfaqEZ1XUHOSYJQR1IGjm9s9QFtkcNJgFMJPEI6bIiMNwIf
HbYRU4ltg9mjjpl/wjl2fejBXVjgFF5LEQtaNLjwOQNTprpWvj/Un74xDDp5hQJ2vNqF0vOihWz6
Ii0zIJLvVavIe0f6qi6hXL7hdqxSo3+qeleJ6jjC6Dv3GriOW8lq9KLRd8Vz2zGFbi9zAdmis+8e
C3UTftgc65X7UMleEPXB1Tvlozh9NKz9ZnCibF1WeQKvIJ5ZiK/UcPcrScFmBKJomglhM7eRwbSa
RY5E1QDpubs0btXcMz0KyHmJCQreKBzs7C52RcLjnGsBUBCXAMwuluvjXeZ7DKCcfryBt53B86BW
gM78nVuPjSO/qklunEMvNsWTHRr5+YpCHDdNv1BlqzivoMpMNRlrIFeqTGddmVWjnFeoeee8P3Mx
39kNQDCrt9HjpbnwpV8AKwyJUFKN5N4AP9x/oyQP1Ny7NM0TQ7ycH0+7zgJtCJkSzLccvx1KDFIQ
PnSESeTIi6n2mM2beLbOpynehTcHSFLM7illUM0uoHDAcAL96pLqKpZ7ux6UuFJRDKcUy6BPkImM
OI3Md64oCguuHphzZA/llGXKMNRrnK6+paYMUxeqO2KAbzuncz5V6tJL35H01GiQeBLXrY+K9gul
ieegM4MUAPZSC48IjpNsS/PbOiCcwKASFadGObMkvP9aCb5+ZeQ7YnPvYgnOy3zWQpkVEHfOFHAP
OpxPXJoHuSYmWx/H8y2dzWV0KPyHtyfiYGpG3p5SCwLQ1Yn5TVmi539JJ5gsjKs4437/9VA95EtI
yTPBUazZS8J3P4I7SvBMTRNvc+OGxMBneDhZEnv2VAVvoj/kQrUszguPz1EcNSX7sh5QpjaKdIzK
yKymqF6q9nWevvnw2D6L46wniKMbwF86DNyqYLImcTUPWrOhffzguxubWrb1yffgLFL0XMmV/sFv
6KV7hQJLIqGzGbqLZtWwYFIb2uxmE/aPh5s2qL9396q0JFTG+al4gv33tmE+bcCtIMf1Ss9ICnB5
oBowzCnj95poRHXHZy/cYK/f2mKToe/5uyxaqZT69sI2hweDnVeH/WG5YZL+z5Grkz/2I6wYoJSi
wTfhE6e9bwzHk2babyp0D7jta9DFofV7tOVZJLmSFGsGzio6peFPr8sdwUkWgXol990UjLwzaeq+
2zs0+BNArWpfUiPofkVX4A6DKl7R9mZKbRQek8uKy8xBCcALDLiQaAVMUx4zVJTLNEVkUE2lbDSJ
oKsYkEJzsx628rp64rIokwqANlqX7+cjWnmWYOJ9WRT33Mct8bTxbBkf9cNVcWiMJr3DsUNHMcHT
Fi0THh5LCkIv/a8ChDP6x5s7DRv7DdqFgm5zXT07AEW4l+/dsaAJijUHFHktD9mOxdL1woB0C0LO
0GpqM2F3bXsYpQGaN04PQfP0vJUYkeoIP/zzyIkbT80uN1WZ7I0sw84bjMk12ypLKCS0zVVewrJC
TBwhnEidKXDaqprgNDOgKs1G9oabIdo6D22ioBA7PhirvLOgkpDQgoLOmP87i6Tv4LDqbW8Aafj2
vjvR+JgQdfqV0aJ9471SECHh9SIKk+JI/+RTMIHPQxNsrQsn84aeRlPX357s6fuQca6HHiTdBew0
UhRqM29Mw80lw/i5Mwsa8beWYk+cBsP+S41kwp1pCAJjJuHHPrAxPkQbSB4MNWlmWty1fAskz73h
YFc7IUzvsPLGDeDsLb94hbyqbLuig+blXjZ4vtXZ0DKpe8lItQlenih4IcPces8qAi0sPanhru8M
k6hVsrt2pW5Id+EIxi63SE2nV5oN59rYlDHivfUYhlAVFfpTvGn6NkGXEYz64LnuJPuWXpcpZvwv
XHt10LTH0S6BJpa27KkmtmEutHUR/pFs8Z4T8t2arQcuwauNdFJWadLyvXWha8ch0tknXZVoUhnq
dRnLBwfH1RGlIhhcGhcTa4K0GaSplRfJEi6T0zP6Jxll6IArl1EDK5qAdL7zOfHxSFYztZRiccFn
A/q8I+v5KV9WeJwOtexPumEd9x5yQvcfq/P6vAnXG5p3VLnVDq46atQshdH1IOGRv9sQ+fvw0+sA
4kRihhDbsJePwXX1Jsp2eSisDSBC+ggS12kB6A1sHdO4PR/6R45jKthPCRdwE/6MkTggjZe/Dd2p
xZzLsUm5c++HPY9hS+ORYZSBnKJc+kGlqIu51WMfWBUnFUYdJJcsK34+0zFRJgAQAVs6iUghtxbB
b2ca9ZFQEl+Xev3BOFK4kLLSr9PtzhyCqYQ9dFClK4X97QytCOEwYUY4guNKfsYku8/nDA7Tsi5T
AppJXAtvrUEbH6sPWoSqMbAMgRamX8Xp6HN0vbpFkx5aX7IhTvx4J7IPPBc+iZY9OKVT78O1LA0x
zzLjjQlFcQH/mmACXnXuIKG+jPGUXG4yEAfAYvppQYbBssHPcJJQAIZEBLmLb4kpuxpAtD+RWsP3
2EN1QDR+4a1Sjnmk4C6ixewVQxdZ6KEGBCK2ZLLBpVfTqmVSWkkHmn9zcMrqUyJof+VT3DabGu6O
uaibap6uuX5K5kIQEfhsCRZHl7foG3w+BSotiRp+ViVNj1gL1FTwgqvZyYKstJdcFXUsSfS6S2m5
NBJL03ToRfRqDBdzkpLuf6oo8DTW9dy3yrjiHIEkxfgx7x2xyBPnPnGJ9HpNCtdVhkXIbpiNeYyS
YmgxltK8VYLWfO5A/1QIhlfvV1YsvfzG9eURS36LbHH8BURv+pS8YKPyPr0j5xfXpG9J7uqhb99K
uspJSBy8r4ntkZ/8gsASNTkxjYIs5WURTa03vjHhIX5LngprqFe0Co5oqC4b9ahqcL3ZcvgqdrR3
hoKRllfC//nU5rmvYSMgPmtGVexJBVI3qaNTYsmakC6Qjyq6LFcWIPp/hyz/KlNvxqCfhuvlFkw3
LAgKInVIF6H/waTopDL0YnQK5g3y/i8NK3YVLD+GnTVAMCbEbtoLJDobt6C8PjSlCyQnvHjEgwwj
L0P2QZ33DEbLnwuYLa3esMYtXcZ0VJyqMc4qSyFhPCI25w9zZ9Jw8xv+ps4C0FkxcIliuJwB8goB
DmBCG2na3WjO90nx6gfYIVTOlAxOjLANgacVe1gs1oDSG3JD+DYYuOs+VhI6sd4CWV/Gx/9b1Lie
USZ2N4rgRJG8JANZWOL0zkhvKJNq77HYOBEihGD9SDAipiCzSxSHkibzcCwEQfkJN0jxt3/xJslJ
gY8euFrsVyEcEWIvBwOnTXoW/BAXDYfwPV24VlMAYdgPdJl9uh5mAuygsggfUrWxNCw5dMDS0+5G
yVlTa8Hrz4qBlcitQVROcoM8V5rmtGNXk6BSK4JZWPN8MeMVlQ33I3DwRnJGvdEua69b4wR00mq7
3zOfNN4UHSyLF/okszeAROQkkJ5IhbZSDZ6hNiwIT3ED0a5+4/kMMpT2MkZJRJ12fqGEUbwLyoao
mOuQ3Vq3NKtdsZwRkwR42P4H5PRKhnMrejABBsEOjPM0pOmgz4nJ3ajs6apghgVwKld80lAN38ON
hkTp4oCay42EnT6ykg5LFS+flEKK2Vlg7AsGaTCH6wZJO8Szv+WBcySqSlnMIKA7byIL8tWbyTHe
9E6rhYOZpYzzka5tKSO52eDLyB9mzP/AP40P6frhLMld6bm3Igz1Yz5WtElDet7CLPKS2+Jt4mn/
TpXqaKyh2Sr0YXyeELIdY0+RWTGVijcbitZw6pP4xX3BtNm/eCW72zcCsuk6E6pzggFYVds2Toi3
PcrPJGrcsgBxEUEuBi/Gn6iFFsHKXnhVK0+kX9j9WR3jur3eEVoVlSIIsg3q29RJV9vl0Fm80Mi9
CyZUjPQRtvwpcDLXxH06oXie3y8LZsgAPWI+FZRypLEx76TXRnSPOXxYmCVDafoZMFW4Koa08qqO
2qw7Db0TeQHfTzUHAjSNHAph8hyhQKx5ulqSIAdurv/A5KAxQo3i7d0U2xbMrBDQVj4QVeCfmPS9
YvUYW8Ou4GPTgqaUu5svLncT/TWgshSd5MVVGCBNoXs4v9nTGzbsclKPp6OgOdoMidh7z+jfD1y6
EkU9FCSgBUeiHWUtUAQdeXrbhvUws+nJh7MC/p0VEVvB5u1eu4ABqOLfDk441Lv3pqh9r893aTFg
t+b7yv58RNAM5LUI4LZ6mDlVVCUCKaloUBUz37QqXsImzphyXnTxluDIZ7s3EkZbVbqR8vo7jnrV
Nyebd0KCxcZK9Q5A6T8eG2GndN+1wY2yDVUncuC68pT2rV5L2wopx2knDDIc6yC/WeQEw/35Iwii
D7TlsSoORzFPT0G6/gmq7BBybIxQFyAwIv/DcAaNuGkI5QyMBerdTcuQK6u7UVn02fr//EiG3FU4
91bflPOeHpF0lf8Jmx+qKfV7CApQIfJEjhP1DfJFtB8QGqSNG1kkqt4VYCoWBmfktmu4e3+qa/CF
Fa447p78BY0IiJPx5pIkrTIno4AQwcXiSzNmutIeDaqkMyBJCFTo9q5GTRI3W4tPaBNSqSndfPkF
AdOg9CfsJwcl0YSJU75zqB+FvOpbnpN7uDyISZbCsbhP5B5jjwfVpDOJNXOSV3Mb4WK6+botKB5W
OjXTwaMd3tC2cHeB8EeAT/cvRfEVnzVsb01AtrJNOiPYYC0DynDy6/p/m4yCjUOShfu1Wl04cxG2
lUDX7BHK1cRAfg/DuGAvQ4HdbIqikuiHBib8OHpqj1miI26qh3pnd6A6BMXQuzJrCH2tlUMJeRwJ
yFfr6aXLGOyxLxtvlPaqymecI9fq2rYb66Q4u94saW5+hn7bRAe2wI5PfVTxQPJuM7R8oW3Rm/P4
8zFzuNxhMHcsMmaC2OmuZm2qnBc/of3bqfRqDQLV+ZomytNLhzclmfyGIuNJ6QmlDByHwJhCjAXd
rTt+RpdM9fenj7wGJ5nebuYOGTlhdL3oIjFjCycU8PdZc/GVrB+NOuTuaSleY/qlUk3D+Jmwbbz9
AP3cd+qo13VM6vwXUdV21AWOO9cogO/hup9gUiQYb4DkcRHiP8RCok0GvuWimHN/lpnc47NfuYLq
y9+hdvryC7P7uoyK9ODxVA+BNHaSme9pjGaWEkK3XEHefFFadx+OMXYXVRp7U1Ux3ctDCNEpmAf/
U5wQLXQEdKbhMiWifmAA8sZsX8K/Q4ujxqRILouq1Mkvob1gAe84Jf+DtKUHFlZS+8sALvcsOdeZ
ebljTeJAH3QoFi5gXnytD1SvOdwDpnFvYP2n+3+BlrGkqqsAUsJ4aZrp7xFl1KxwR5Tn77yl7R5C
ZYoknK+RpHv2QWaam1nEuhtQ4HQ9bJGQWC3bJvmGwMGcDtvduq5l57y5f2qB0PPIcIAL7dLi1nGd
OfTsRHEHH6pO1ikZAS9XqMdQNgKcqbotIhEWsj00P40BFkalzymMOdJ5fmaOkFo1hK7Ooup0EX47
vNjuMhV+cL/v6StRey4PtM2kIRS4G9GK/aYEBGgKw5hmkfWV1jqHPWpveGuwcDJndIn4oPMWKI82
7BjOix325+h+NoA+82P4pUtI1RCm/Z58v3YLts0O4waKHnC2Pnvte8FnwvSfoxNzWibS9khttMVg
eFmhqHme9YR0fMf01eeVBjHbql1moSQFd+xLGfbXCu3LRJ6e6G2gFNQpr2sPzbOd4v+XcrGH1ouc
FsWuqMWIxOUw0eDQjguu3qaEQQ9Q4L826MNp+8O/v9b5bFMD3jPZE+KkoOZpLdRwqIqXSTBsLDCV
N3mYOTQlJ0qWv2O3NjZonPKUx4nwLOHpGgBE0ZhYvhtuVa1fEhzs28+FeCqpiQKc+j7o+q3ug9at
DptlHBbcWqcFfwaNJ/oRkzXvrgJjGUeoAoibq1U4a2P4ZTvdWcWI3uRscALkLHarJY5CUtPb9yyB
6PD2M5uI1WZQU4rY9329IC233H3BMyeYfiul6BnZJZGjJRHUgaY3+30pg9m62t5D8rVlXk5KWFuB
VTVrqTIUyxYMghFZl8wasMdczJdWpgy3RF8jQwvaH5QlrEWOFYBxhj0oUA+pS3v0frdeE/FgR0XA
CqXFmoLUCtWP0y6o3VndpR0846jxmjwmR4lrWlmF1Qkq8SDs+et/FFA2MUYn7HBbUQObVDzuxmv2
zY6OBt7OSRB4orgcnjACbZEZNmAA5dqxJIFtRyyG7GY6QznlEriDI+WqWkGIw9Gu5RKst1rwOyRA
CtIziqw2J98RsDGOYTAGjyjlYelqXEvMcd5o6Y01W/0AyrETYdp2jW8V+njGdKeKU7p/pRuRPMf3
Bmdlj6Y8SF9yBzH3qcEliYj54WgOZiQnWZgwgrS8G8eaPgndrU0m3XG6A3U2pC+zR+cniawjl1T7
W26020phfZ/7d1gUhcuooU4YUzF9esDkxqvycnpNCM9p1/MDtu1dzefC4of5dGvzc3GrmjfRyRWS
6NPe2ktUkf/e/OoJQmN0hS38dz4bsiREyUhoK5hbKF/mHkfKtu2rYd73lzbnbHIpq13I0q12NRfi
avj3zzD00HfAz0mF28SHIM4vqFBRQXY6QpV67BofByMz/4/NETiTEklx/oyJymHxft+GITCjsknD
P3mIiWnk/Tow8g4TAzgCgvcbEEinhR3v5giZt7Tybhvi0nwelDXlAGwLaV7414yJya8XEgn3wixB
u7ujg9ZUqnVXf3eMpiXE8u/l1gUa76ukOvPztmfazm9Uv67eQIZ+hqOMv3LAnK9CNgcXz29+X6DT
kg6GReszPyNS6Be59h/xYj5kiGMupX/lfLfS5QHqgHFNdRsxUfKWnVZVRLTgJwhyWqhOARl3ozgV
WXXPWT4nLy07aOM7rohvpj7tERxQjnwDDBjl3UJWzXL9ITyC3dHhTvQcW3uHlEora6GrlyMqSk5C
cPIKHr2+MfKFE6PMWN76+BnS10i5mwgeiwXJ9CumNCOIJ+7UE5me1AYLXX3MfEOvZfgXVdBMiyHd
nNnao4MOfVYa5d0LYQPYhCl++TlSwBd97Nl0AvCuhfEi6j95N47YubOOyr7IzUKZyiE0E6On3A2h
9aJynE8DZ2DGrCGLSwuMTVRw6Cq8KatZVZPFZrf8gIh6TTuKxBWADxk575Mg5tXyr0nXfD7Zb3yN
5wkKmhGbOQjSWu1MgO/UfHVcV1D4Q+yv8Xh+CsSis1dNTjOdaBLV6ybJU9Py5jUdILyqncvK48dp
p+MTARstGz7U6LlrPUXXXp2AEijs5OakP00cmmbB2YmxpzmnqOkWvogBmuZPZbHw6ERHo56I54Z9
75ri9nVTVoIoU0NHhp2cBo9fbO0eq1dvs3qLmvPS87TFVrnHuuqiVNvMLO6jHKNpGCKmcODQlM+r
IZ2xn2KVxAUVYguRZFyJt0Yp1IJacEFEqgNgfVfEGW8okN8zFSqOZLLCUjeRiAjzk3ZvNCUQ7962
B56IJ6g8+kfYcaeqHQ9ktIpNiJIrSBuDjeGyzHwkMeuGrrmeTO+LxDnjApiEbfgr0T73fhaGrPya
4299o03v2yvfnr+Z3hUYkLofyVR9pI6gtVoUZfDls4B/QlfeUvsdUa8xkllaaK/vGzS2wfhnMS62
IDyXU1tv2xC7M3trnq3lGOkrz0ZcMzNye9DmO2Oemd7K7jvHfQ7ZeUT0Ir2qS5z3FgzgrEZNL46L
7Kl7PJOzlf5emnbCLBhmXcmpTSLkMaQ0+bMw7St1cxfiR6GzHBv2wOkwv8wlFWUIrt0tHHiS7zAa
uOp+Jn/43nqaiEC1wxEjRVfwf3U2prSBZDaPUpvwiJx602NT1N/eH7YDQFkJKAsAfJ68vl47J7wx
BkRzj7/ii9atd4uimkjdjyluXNBev+ZvuoN5Ve+Cw8J2XIfntra3/d+IHorvDJN6DoigM01X8H6G
BkfE/yOJZO11lYQrjYDbqCJHiD9WbPlB0ceLDB1sqwSX4kft8iBE37YBGtDMudzxglfFM1V6czcy
GUhScgCcZY35p9MfOGDX0EfB3Nvn/+B/1Z8eFsIViANp3nYQ6qmrqsFu+bsRLDYUUjIXO5sniNkS
sWLpL+64dWJXRYZhcpvSFw5y7IPUlHZNWvsUMfibGKueceMSZ7/Z6ZWtUrluEGPjUWKuUgZdoUHj
bzoQeMy+VxmKBqgqtf3EdmfEx36VgjQdPTKG6R1ctQWNg3EnNg0+2eoCha43FTqWJRJKpexsv2+M
mvctfAxqdr6/7vS/7xUiVw7wBB42KYdKdZfTkWrplN9s2pr99N0Ad4V0SEpPF0Axdm+letaTscDp
BZ7zXxRKeqhT0u2+IwjAu2TYS7trqfsss9PJKKVXWh+wr1/DXK8DjwuKBMaIhF4evOoUGzstwmdd
z7iL29vWpDi4rZott88WNrqSktFNe0EoB1EhnPggntT0BPkgVBq29XmVpAb/PN+kDLVmN8XpRhh4
LmFyQ5lNQhyX18nhQWSh/jYxPT1zzaqIBLCUVCDZR1YEXUiLr35xZCwuBA5SYaGVgRfW8uQKujrR
zZBAQBDS9NTNbbVJ74NYG/nHtuEnLbbwJKF5oZ9D3luKj/Oz5G0mV73zLkeZfCvZ/9jCHG21RlWF
+1xadEUlvgvqQBOQAxfJvxK3xJ0ynvI+vswMFnkbgWApYgBStd0qMFNUzCwpE5hclVCKjHQbkYab
k5bKOgLwZdvGxQ1tw41+7gm+RMUAdL8E8yx5PUmh41hRMUeQ98amQqIvjzvg/9SjbjUEny8vXDCM
sZQkklD2I3+cGg7EZNuy7Hpn+0x3QSbpxm9lVD/GtV8qk8PYh4zZ6MOIM7QBiQlTmKImdYw8zYux
m4pzovXMexni/FOvi/i93J9kWKywhwrE59gmqsCRnELbHEaib1MHRBsxM/BiIsqnPT/U1kEYfdnc
SH039cJcK6YKC59PJIpyDUrJVeJGYrEk/7cBJw6K+70nGjpLxihkwsN2kW8YSK2SzvVwlWT0owz6
2MvyNELEYiqI58rxVa/stGCRiQwYN6e/ad6Csg6scG80TyADzdXK0veWRxN06ZE98JiunNiuirri
mkHR9440w87ceITI5l6n91LG9WaEcsBHyP+sPnor6x4PLzKvtaJ14J2OxQ+coYw5EH2MFPsrjJlL
2r4v8ksoiLR2MQJIuK7c5Plkzuuj11s95Lxgo7ez2Wrgrhb7NyKrIyWEs4Gfk/4kujrcYS2mBjIU
c1ONNht3sEv+0H9JqaBiB2FuuYJRMmbIHq37Q+tYt1hMxIG+dMYNchAmfmROighfFjJC+fkiD7zY
n/RNDPceoaRI59ABnBVhC10ymE7dBkKVA2mkaGMzTbCU3ubt2d+4CccCRA+7gYQ9mkrTYmaVHJne
A0XN3NmnFSMoM+qA0LlVebkZ3/ETNfctK8OSmLPNp6sbSVfRjdrnVFYHXhxJYOvfVUfe0KJZ8Jm9
Hwpz9AbpkK1Ec9G5q3F8uv8kr7DFhF/5YGk24T8USjhf9SluZ37Ug8rCK6CugnA6GTXm+RCqnMxP
V8jo3EYleZ4q9UJ1UNjh/Nye2x7cHmMks0YkyTiJ3tFhwhGwGVQW6WARU20xkGh53bE2PPogn237
bl5x37syRg3o17dyUs1Hlq5+9DKWOmBOYQ7UhERrBDkjAIB39937K9YrXmjvfxPUQeFG/j3lwNgv
mFUoOPSSeSM5RAHUbHgRZtHyHqB80wACkCzq0cDkDK4hDAmo32sOvC5eu79ccQ8yEmDRk9wh4RRR
9eTa4Ad0XpaGSjdBAFdrCAXIebRiaJDoqedt03o10dDAlg7PKfJl94rM8+a3+AFr9bZaq9gxPOsb
NgG8IWHfUAd3EW9x9KoLNDufgsvZaTUGf7d7Rax5ZMbJttK/NeCxrZnNDC/umEQ+yxzNibDhidAn
AM+kttulmDCXve6dQ0wEQPA/IOqHir07OxvQvc0LEhisI1PO+VzguQGED2BztrzRjvnvNUNEOjpA
yUyCrgmkapfzF8Qs1QEePSI/3U1/042BL14drt8Lkjc1EIkLi3kl2k8SljgQJu07G5FVLMpGrYF+
hx0MwHqFTB1zJp9ItWaikujLl3WCBORJsbO1oBw4SAVoWt6unxfPEVCXoLVcLTw/dNJfPR5J6SlR
DYmZBaGMO2gRbsViOxKWQdRj2B27JjWVlMR4F4/5hMZA3sWR0RQa7CliHgQJselbtuZwMcmYN4IN
kxIOyK6QHXkg0Y3DEWQfcmpXl6uXbrzX1dwspRdHzaizI9b4gV4dsTXMjtBtfc92i8PLb+CkXd/B
IT7Iz4OdH3Otu2PQqDSHkcQog0No/H1SCBieAaiWVlkTX/9E9st0QF1apL+wZLbVSwQgJQbHDdeT
soxSSDcKuPZyZOrID2BuTf/6lpa01UD9G+rwbbjihJM33H4jceXqgIOuPImz9N/NxEp4s9+H3fSY
SzhPTqm/bzEqlRJjiMRj0SjtH6PSyXtBNs/EvNIyYhtC2X5jxlDCTyw3HxdIYfVqi+lpLRCbsEXc
ym7INEoNjXHm56QBq7ouk6+qRmZ+rt/glcbVpC2VKRObJ0U2FDwpI5zd3HrKDzJhXyzhkL9yKyVk
F88mM6qEy4L8tP0iugii5P0LT8nzaEusPV/PlMIiiDI5PF28sgF0C+8WIzVQaOY5038z6FSJNJeg
wIx0JXutYdw5Vdmeu6EtM1aRFwec9oa90zqoK7Ty+WnIiAFaeD3+cNay/6qFhhYuFz4SlrybvrzZ
xt2C8nAn1XR8GobV7GuCD8VKST7N6EzZ6bL1eXGhYq69FJhuWpDvUAWdo9FsiemE2KpPCpvNGt5U
/szJDy6rWcMa4QtE1sKE3QJJVmMrGUP94W5JO+C8ZVdnAoQAjYWzZEGhhEgi6QRIVDsM6g0rPUJ5
owrXEtvkx8v/DnvvGO3b4Gafplo7DVQ8//wOuxZMgaMi6XQRY8n7glw14z2l5If3oOmOAOF7T3zC
s5TLMpPFd92JFuD0HS6dVmotaCdwqXaizl0O0ROuPNpVqWQkKqdL9H3igcn6G9OZizzG0sswViwV
ieE0VpW9xHZetGxmGdtAl2wV6f7A2cEyUZtOnpW6r/dsfEn/bm5iP/nxWbKdJBq36NWJQtxBhi4I
/Bl7cIGjlR4e8IzeMeOF9PUUeQo1rIWEbZcyKYV+KJidCDDOfbA+TdhPQ0RAmADkbLpTlXNGY/aL
2wjkZWj4m9VWj6BGbO/F+QATPLauuXqrIOTkX0fteKVm5tgcIz2rf6z7yAruDCy883i+LR3j2z+9
wUZPiMvFKgSzMR7Gcryl1Yj8hQSFnwOjCmCnQggnStdk1O2uxLIC3MO7O6T6X1h1SUcNzPPfbC17
dcBBPCdSYDN+Od3HYGPeUhrknRRFGkzzKtJ9nTyHN9SE0UX844Sb3uBiKjxHndlmIHhKLCzhqgwk
zZah8aDuPbWBLMgA1dWMDegcr2wbhS+SuxRlSCQqapdHFaATWJtQ8l6D4WCWVG4qBAkStHyPqmfz
Zqn1tVKsI7/bBioEGfWAk+YhnsaVV7VRaA8pWX9ylsuRrgJ6gcJX0ZA+C4mvCyH7jdqis+zSnsua
NpAEaYr4ldx0wc+N24TUzvifFgAkF8egDFDYfuZWr58aYqhTi90OliJsfUEcbOpmG6q57rs1SzzP
SOknhYCUQSj2F93vrRBCCOplNoE2dof8OsUjCMxYNtJajyEShJOJOVd8fQnxIhRUzrS+4jCXfZCv
oFshCRYASHaTcEHv2YYQY2fqgogiC3NMxqTMMzffghRxqYkWep2vJ8s1RvBjbsBPLDcd1zUzoByG
B3o2mSBAAAfUUpEQn+c4/yMN6BxrgqrLmOEJIXX5i9SoN9qBOEPlN4kIPJWnTQXumTjrWYXTCApw
QNCWjQyGeUvlnHdYwtfS+EZB3cDi8Um71f0wna3DD9CgmFJC5aAhP563vPXiwSKiC7qKJLPkyPDc
N/XQ4vG9OjThs07BkXqdpxXzxpbn7AMMPvzDuZw9AowAawTquj5jnchYzDydWHuXJommdODsUHwc
5UANcF+Boed7sbOLSK12n+qgseHJm/mXEa6Asju7T2B4FIzJQ2K1FhrvnXm3zZH6bptczBbk/uOW
AdmKfw6gFCbh0s9q85LweBHlZB9maiCMdWR/flWiT+Xsa3TIY2MHoht0bD6QEktAYSOd6ZGGNOmR
OsOpIy0j4J/eSYGS4iW959pTjWRdxjmXXoCReXWZieAlO+3cwG4AxTN99YspjKx3EmwlfIAG7xDQ
nQ8LhD9P5/C+RsLKf/xqKb31bV0VIPq0aCM+F6URVFe5wSo0T9jiHt3337yY5+Dsi3cnuPSojA+H
rCJV837HXacqLeMeNlG255uItD/nKg6nW7WS/kvH4xqu8rjdx1tHX2oIE6w52Q3qwJHfGuGmlfba
wg4GLRZxTZrMBAKw3ReEYyZUSKbplIofQnCivSscQzq3T+SwJOaISHWu6Ff2ozIvKjyXdoyMjzr4
SXOXe82E/gUITQ6wBvlhU2ZB1dxxW3IS0RtNP5MLiEERSdZ1wTcDWnt30bpy7VAbxYBfQe816K/u
BsExzlwhpyRjDjPjF/p6giCCQCSj4wKTwS+u6TavjQEQSB2Lcr106t1wxruD8zoYRgTVKQc5CvAa
G+p0fSzVCpe6qsRljQmZ9ma6pbmz+yaLcwizw489q8JIWLEdik3oQLGPyruq2tfkPAL2ZBCqo56G
+8i7QdkeqHCPQD6d2NViIyFjrX5VdylzVaGqDvBcvDu5FXezN4SfcjUN2yfIM6i9c1sLnYzMjNr8
TpDfqfLUYMO4pS1KpfmZSbHJ4GW6NRBPik0MWGS8Uf9NmVQOiv+GxBoQ+6I985QOuoX5odOOg9n8
buho+/7GQRN+CcZ+YwxO8IzEKDm0AUA0tOfpI5BXEVBU9MUYtxUOTxmwePQd41zGwwAsPDXnejCL
o303GV6/Xvfc2pwUN9vq/4rPCmnEXoo6IE6rqwUkpR7ADtevVjT8ju4SjgAt+nepmjA45UvxhV4M
N70D0/0hA0uTQt9Mf1/JcaPovYnHdLN1FXbfE5lCBjt8zrzgx9VkZyargSQjt6r7wVbgLqIeDCK1
YihFQLEnhjZmQJDymwFkGJHDSL9w5qP8gg6HfUa3sb3ozuUElBeJ0ylinBBnCe6SL3gZCecbxlii
ZqyZOrz/SNBpQ3FptLTcoSgYWHiPjIk+SpF8MstoNKEYQfItuKorVJDAnJHShVGrbm0wq65/yY1R
5f8aptdpnHGI5akrtlj3+8fSWdqi3vA7yjEgiDchwlx5RA9UyPlZw6SKVXq4q5QD//SV6XMTFXfS
qAvU35fD8J/zrNglPqQ5JzqgKbXB8CoEUngOy678+zhafRGx+8HLohuVNlBIWK9dJWzDNdMAZ7Ax
qPsl6hsKsmL9N+qh7W/ND3kNFuo3/chGbVX0thmuHJd9ETfVcPGyLdsGSfGXZQKmAGue2Eyn++JM
T9eVwJLJVxIRi/EZaMNJ3Rxa7/In3dgfPI5WACTofEEpmex1cg3Vnxwk8SvklQFH08bcgxbBoGd8
9x0e8MUGYohmNjMgUcoEmerZ5A7zqvSnxsb3I9DEen6e9VB7e0xh6OHvEbgprnJQYwR7l1cUbA1X
YHj+x2QAUWsm6yxfseN/GhZa8fiX79tPHhBBF80LtjEyFyeXHPI/bpBVQiIaCJ2gBQOoTs66tV9x
FHtsd2B39MT8kUYlEDFfmttqftAgeuqDfVDbUD51rIKJEL0dWJIgz8T04/pCcQX+K9O0yusI2uRv
6/YF3IuQB2RU5A+ZckfPWUumCAitaOGVuHIuaUoNryGpjuw7NnRIy0pCSqppE/Hx+cAOFm15PhGg
mxqJ/n7QZiglqKuBEcuCY6RxftD7tSeyWZF/+6eoriowsg6RfVYBVT+XEE2UmisT5srK28rO+o9t
/FHq0xGJZhYQsWLOBWki/m0nkOPMf1s4eJvqG6mNg4q/cLf2sbs7ETYBkjBvryn4KS1Qk8X3jtYF
BQUI0gaJo/2Bfrdy56p1zueIrBPCEte1zc7z1DcAIkLeRfAJyV5VPNeYoJbfvD96un2rWBFcB1fS
q5O7jMrgZI+HjOjORka1tqof5RBoyOjWMo7xJAqNgh7lA4df7YJF1olo3vQg7+znsVDcosZuy0LP
lsn6DCc8Gpe04iWEsgHH2yZi4URPtYInzA3Zd/cWdX2MjNSN0ISjoMcy1o5aGFtPK8aLwA2wazXV
lNyi4eJsIL0NZG8KmJhE0WYz/42ifgyjTFTkSpTXY37m/FchH4RHWR7VmkEDyc1rEYvtR4OVNQ2a
DKINcqjjxqQ6emJz1Laf9PHngn9pO6FuVN1SEbzV7aH5ROwsykWsbFVmxr+K10GV7s51JMb2X2b+
0w13QROiJNymgSVgftnAQ9gH1V0EV+pKpG5CIgujVVoDIHr0b8cXG5WcsKKyvwSWwCeNW0bRP2QT
cq+mnLu1pzVyvHgRTZtV+00ZLhjyQRcSG17FrAlw5r3Y1TsjucdhzG2//BlRnj4q6s129zKraoJg
dEpRT666Ucu1fmGEeE+f40pCeFCtlEgnaePfZZ20QVkVj5yQEPHUK3htEThkxE1YdOFnx2gUBznR
dhLFwvadW2g6vBVd2O3265COK1LWkQFNm7GLjjoC6MZCi/kQqdEGJmirFdWfcWhafNve28q8MhxE
HnxXqMaV7p0/ckbmBI6FL16aPEp5ON7Y3J1ots/08H800re7FHBQ8mQ8jmD/u+bvRKE5yKg+5v9h
iS+aiWSAWlfEQgEU5aR0tnMpeLEfwTaNW0Q3z4fCeGxNtxZBO60Ihvps6AKyEwC7Y5Vr3nvwvWy6
9obUHwZS8OMZb9DFuh6iLhbC+5so4/eblN9d3VZf9OlD2QulGCFkmCseWJVS2d1woPYf6jBGxLH4
KK1fgSsYhRNper9R0NztDN1rbyoI+LBQyaCkuLfOw8AFehaiZcuF4WdHJAHNFiarsgXVGrgQzgou
14SlqNEdGnGbtjoDwie+ryGJHuO3X7RnrVrOBFNfW6wIFi4LXs7boj6sSF8FY3krEKmK6XN9MXtt
EgsBn3O5AHF6gGjbLyUzEK8/CA59GWMBA6YYCo2g3BLcLvBm5uvszc4tlSQ2yX1fBZsbmfeXvbMV
sOKFaTgjsBzBksJaO7WHgO8K6oXmZyeQGLjFpIHHvQ7txM9ErOonwChOmMt+O5l7xt4HbpcEDcMP
K1MTOVFhrj1WyYBsvDmledJz+w6dSQZcAN8iouYL02Glh4Mm0CuNl+Tgjy+crsFimVXJ9pNt0N94
qbI5o93bc3B0YqJsvQSyFxfL9JjXTgN3saQZqyLIY61K4AiYt1p1zYGm9FmDtVLB2URtPAZbgc2r
ErqDYFnDUiLe63NZmcZ/5BXQw8oS24G4+zoFt7NxoI/W0oig7bBoCgFP7e7FEqcmmIpro1mqpj7q
ocz4DbgWTL/pGhmwCuDY7LA7dyhv2Yh69lKpThRLB3Px3dJen0soN1be+g7amIaZs27HY8fotZJu
KL33myFP2fpIfiuRmKJegEFOKMWgScoivhzgoszEtkA1cfx71uRTMVskNOieMJ43u1P9ZP0tYlvS
JLzt03bxPfYq6GTGAkL8ZS4qatitm07qxzaPE7Y1BHMUsKGAlu9bNPL7+HAx7IUcs/2KSeIe4wsz
TnvS0sfrbWLwNziqesR58d7MleblzU/zUTZywDFJAj2dGhkFBENe6CTW+IPqs1wkabvGNkvUo7nj
CMQPsQ/YO1ii8wTWB7FpEVI6bsAqnuTr3SnWZLmdN7mQLuE7gBw75S8CoTPpWLrEa13udAL201Ql
onCVDjQo9JHnre8iyBd1ss4hOVZ8GbohlLIm8vHLZBLbOH4inI/kI1GRosW9/p+cCABrWhVqbp9r
o9ndlFaChrHOAwK3CcMkStefBYZM+7SS3oPPbdxMLNS4T4qJXVJLFNTsSwELVVcTZ4y1gC/rapmz
Pu3SfVUpH5xRkduSP+YSEwxU+1/6yw5M5ETgFDOz/C2iO4zwSrmeUGgRiK71/wca8njqDMi3K3GH
QbHY0cluPmua1R/MHdD8El21YClPFioAHNzGXs/OzjXpFSDrLkbfjIpysL1cQ9aHO9Tsvh0KQPJ0
tNym7RdNbGsvVkHJRUIBWJqLS9Z4TeaclDWzfLOVmpTzCMymPFznHE6IM/WFvyGsKxkK2BVJLeUu
RplBSKPYvf1e8Dq+M4LTIiHNlAkKZD+pKNahvH1shJdAMEQvxgthuUOAhD05pQz11heO1huwSHCZ
V1fiT6v/WkFz5M7rY7pVR1e0TuThI3Wmx5H+BaflME45cScThkeiChRFhR1BaCbP3H4mrRw73UoK
1HVzwbDRVr9207RgkLSLChvg8eCpoYeA/1TfyU28LDDYzM7hTIDO0Pp3l4UR1B/dHVtS+rCIW/jk
yOeUiJ2kToJLHKNtvXArX6vOON9T7IRtPp1tx4pTIcAvU8rXVlZuv7YRHp+tEgxCgDS5DXxpC6sx
26pN0//KCCo6Rs9nI7hXKo9Kpr4uqKxZo7rPglXRuMDF3SOCjzS1GL212rd0+EdfsVioE6Y3tlSu
2Se2qR6qaz1sjO8hxfpokwi8EGXYN8iCIyfL6CWGjog/NfFIyDoCEgzhyOYh9MqEUWFMIun/G0UI
FDGq6lfAslzyq2O8rkPs9XtQUZwYEq07OMuDJd4Xuehtwwsp6H7SKlPiNCvlqe6K+mR/TFyepgEn
SD3Wgp7Dy5yoaLnRSEdO9rM/PKxCKBnqKE18481A4Dr1SsMofIxRpxqUFx2dgxlKvPijezLwABf8
y3f1Z5Been9VMLS9iMYh2wPHPWJNcbLLI3G7MB7qBl/qSLYenERpmgptKcMT+8ksf7iVcveAWQ1N
s8L4SJXDvzYy9xCA9qxfX5BrpdCTWMlLn1nb8KRpA+KCWL6li/3+IFE2VVqL6z6zrhK0jOqhp00g
0qMH6wA9NqU8Gv5c3ku9Sf6y3EIq4mxDgFFg/GPSolS36fNOYxjIUNmtOFlIfq8qgX68QWBAX5Fo
7KCqoTar79BVS2+709xO1eiOrmjgk1r3dCR3ktxidZ7xhA4GLugTz/KmWKaJB2c8sJBlHg0pyw1L
6xFdTga08Q2B8DKvUdgTJd38uXNIJK4pT83NJRlvtzC/kJO95mZOZZif+WJ00Dcn9ipaenkvoZrW
6nVirJ82ry9gljHh2WPOC2TSMCQ3+ws9xYU8W8TCt9pgb1b0ytX5D8NLU9YP91tRu8xpmVxDKNIg
UsjC9pn3ysz97HwVXpukYV9qCp0KC1EEES/ucLVYVs5A2+u7Dauqur4oBhA6q04i6Ny8TXas8dZj
3PQZF4OGvGqsUHAJkAarkI6mLbkdT2qu4A4qgu1KMiz7z9T8q3H2StvajtVasw9IHfDl2JtgHt5v
EmJtVd2l41RZYulghwWgtTfXRMtf8hexyymQXpFpA/vh/e5Be8JR0HuI7QQzfylb/HbJktIFGO1I
AnfBl4HNdu1gphV3gg+vwrd9i1w7/xer2HmAJVIwXi8L1fTWWH75t40hMNZiortujear/NtpmVs8
4DoSIiTRxBTpiycXGyxmKF992H8lrmHx80U2IN/PM27xZEDPrS4B9h0zAZDt6CIubdPooUsTixz+
zDbPe0wVBfsWNwWbvpO1q4pCWJvvKKQzKsrxD0molZoTprsu5wPFzm8ibVlzdDiO3rX84HvJ1bJH
tJ2cNuhD3MaqG9KHKiHqV2KJ9WiDJR7Daf6BR/gIlI+O2vLeFhYacuebla8O4hrN7oQO2VdMNPOf
6PcbA9qamYAdI2qF0kA6qd2yBc35dbxPtQkW/+cnZ+05NyJr8y/ZAntTQg4LFpkOxjjR6tA1rOJK
GyCXGrDeUejP8OukqGEkCLlurNbJ7AJsJ0gKeQbjmJPh+mHNe2VSP6IGvhOsXKcc82qMoiUbHcmZ
G/F87sSefD8hk0Yrm3fDjbfQbeHvykwfdKn/ODCx57U4LL0IZnljkHgtLRhOCf0h/wNzXzrDNvIf
M5ntRhawCREYnLMEPYrkuMRKeML3HNW/g4vRM2MNLuhikzn+7BMhApNizTDY9O0wDkuRJZNHHLLa
ODxTFj6F6r+FFNDlAGvKaQEWXXgzBLkCAumFyeBKdyHeQvJtReXfT3CnaO9wAplPMwfrUhG/Dv8S
h+RWvoRXIGpi9O5cdQQmpLAiCqB6DItiObJfyPEEXM6wLvkolelOK1EAu30/rgM61sqvP2fiAtB7
daYdNqR5Lqjag7TVPnaSm8HQ3neKmqtV2GXXkT/fqshzi7l5l9tYAdvvHsJCgs8HU1g3UEY+EBmf
Vepi5SIKKAGBsoZShvM1nF5PHBiS0JC8LQkvpXQToJM6/iXte75YmPhQbkrK/GAb/QCM5ENEAPwq
Q7a2jWj6Wr1MClia94dV1ljApy+BWoYSVFMmFWTpOoUY2sDh0ctDzjY0SNTcnMfS3QOSYU1k/D+W
bc6rxkThC3I61sTyGaipg177bP+FxHdhP+mKucRCb50A7ki4lv/jG24a59LjWkkUWiiA/jQVw4gz
FYLOF1SZU07k8Ml3yn3GlSIUjQBh6MIM4rivyOIuorMQaL+XlPFGfxcXBoJKgVEyQFJggwEgsOc4
Fj/a+e9LFhAOkiC+uz3Y4Zo3IxDTOwkuskD4/PMAeuxHFivAMzQUCnEZIonmfGLrWvVmAMVB9Iyv
Crj1Lyx2UHhGTobVN9NwD2XIj8BqL5I6E/K+q2WCNWAWOFo4Bh8JNLNTj1fRM/Tcy5vUhpGUlZo4
MOpwyXaJxfl8+FBu4f5XGJVGDSc/uRsT/VBUvV5aN9BZz/OJd98F3w5CyFFVZY6ZyZjCrTRaPurR
dDdIw9uuI9HpIialn0jkMUnZnOIuvZJYyadD4h5ZDC13C9BeB1ihyv7GYYGYSL9qARo8fru8lwFl
3FVRDp1wAWKT247nlYhfMCyXozp+/7UYW8NhfkRjQ71cQIj8CCByRGhkPX6lMH5L4YImf5lu6uDQ
xoEpIFWQFqR5cY5UNZnDZEiwN1TNMxAgq9FyDcJWLnKmCPfWNzIsbt60BIPKAMNPnFrb5hy8/Upd
+sxpE5ZNy5oWAr2wezSuW8PivXDcwA3qYTwFdPgZDCOqY+2vFRlk+ldDm2KLC9EMXPHh+qrAXR2K
KoEFJbJrAt37/tpwowp/+M+/ugSqcsJcfxZ9KQgvwfETmUQOcGP/4NS4xDLBPQhqKtzUTAvRsijy
fn7yk+0n8SEcN+owVxqAtTkvmv/6/OuwRgd+wYIkO6nSFiauv5epswdQdg4GCNJsvligK79Rpoy4
dWpssl4w38ROJzQ1kiWH/Bzf3+mC5jjx6dVm/HHJ8dzVosZiZCy8FN3kuRLMRE+hWAKvlf8ZXFJe
t+wEqSl0vqa8gxZYPiLPij+pNjVL9P3zwhqrTAYXZ6kKHiCHB7aEVLlUzFoI6f4s5Yq5hWEg+a7/
juDVh9hoIRM/kN1VYzOqeXUI5kS/bcEhh9cdIFgZyW/O7FN7Nvq8JS+Zd9DeB1+BmUOQoCS6hRkG
CUJxma7rge+yJlwmgrsbfqAQ/k5Gufyk4+Vp8/gz+bNytfVRtN53G2/4hixsybaUv8v9MTNpiegx
kciez7iuNw4im5i6V5QjBchib3rVdW/MlcLSWiJbqgQdbDPYZVG1Bn0HrCoicqDBwEp1/aXwSfSo
+D0e69TYQCc0PGNlmHXuAstpk4XWCD8c2GEYB7XM/C/cemQNPTN9njLODShY4CNLEI3pKIajjx5m
C9CW+TJdeazlh4LpUdeMYTPTxHREGnhjSEdp0jIdF/Hj9F3AFZGwZWA8IrxD7tjKN79oPuwG0q9q
FD3+FsQCzrDbP3QytmhS5H5EWHIvhRvrloxPjeqdLggLan2I2YPKYKNscSsMDm7g/b/MallOiIkZ
ce18T78D30kQ94sZ48X8MKXUIxQP6+UzFeG1BeMAsjqyhSjF+cDqRUq4z2HlBFVq7trcuqKBtGBw
78nqIng1vrjau2UWhE1ZKuFGFAHHnC7EvSi57nG31Du3kvN6cqw4VtLXsOIlfa0Uo227zS7jsM1N
0kjy0ZO1A4rk80X+OXu1jwE9oH2ogP6pWOyd5nLnxGWNcxe/ycomaQJvXtyfs5coxeoh/YV6flFm
8sjQnZYAXVBXkZ05dGwHLUVuAE1bdSgML5ePDwGfmW/Of4hB1jbMNpu2ZtByxYx794/9eLd6h+95
5BMHjAwoTRmgIPlit2jwD2X0A8cUSnis8AzaU2LS+e+192XAYVPAj8gJ3B0ZKzgOq6gy4Ulcecog
i5pbioRxQd5U6qvYd3+Ej8N2ztEdiFLpAwIwfl+RbjPTDEf7d+ia0DdelNaEh/zMwSNbWXdC7eIx
bWlPfPlA1xDpMKETYNOBovi513d8qqEGVgBz+3chHm1/QE/794wf7ulSLTAkKeOQG+/7de0/AtT6
Vv3+v1UbZK2OXzRHmes2YMD2EZ5meWzyEoHMcJEmhFAO5CKK8rhLT1Utn6GKdYM14A4Ue6xOav80
AbGon+PdNTsQW063XlIauirNxk5SIaHgi5g8T40mkq3q5myLJuJsPZWIfQPdAt40M1hg2Eltg6A4
GilDDQW7JtLbC5SXPILs/mYv87wXIdEGCvAihbkunckHn5QnPJhylgI41nGNiIqBIUjd5sxz5vX7
lNFRMTXWx2f1YEyGx+NSraq8jO5b4qVYUJQygVk0awWeLP0M0fSTIp0L5RNcbk4xHcksceeuO7Pt
KRrNYpI+GLowrrQWT/nfMkzNDTHwdAT5r0EwqN372d+XmV3PAbMOxYk6J6BEHxo/E1oeazQdV1fc
4v2VvPHO9Bg4a74lYRxsUcJ8fX31hHID9SRYeGhuzYNJtS2BoND4EvsXrROQeHwDskI5bg8K5mz4
O22x7ujfXHgdHRVAsCbTJQhWeBRZWPRtFABmMEr5PXILZKKgD3ifyaQSR2KBxUhgE9dQpN0BWsv3
iQlsnfd8FS0bUmT8k5uGPgnHEhoJr1d6E9NE5dvfezZShqQpAQiaQQn7yXnXv/nMQruTZ1R2n2FC
ZnfpCwrWkzCJN9tYCmMcZ6xXm7jdV8NOIhO+qztqNyGGOXx43J7UNIB3FEY5Md5jE2D6y07XACBd
+D2pgFm7+8b/G7CadY+ScajamVKmEsmZQA2Z/WbYYsEr9ivbJOqTZG0qtcrkKp4eJopCXDqPA7KO
pKdPYsTIeLSd7VvgCbfo+YSPDC82gihPE3nwmVW8hFJZm6K+Va3q+vNMdPlLHLO8kHDyRTnzl78U
mdRjBitX0tPp9tuq6TsP0Sx2B3zwViRxr1kYiHfzIYIIbAeH3NeTsY85v7MaxIKg0phTrthKLYDK
GXr0wpmlu7Vaaa90GhkbPEdvxZlWjdnx6KL36U+FxCw5azLWx6Kl3JFcbpBBl/d30CCRxDPZ4EEE
hZYo/EgyFJydejLM/zZFPm4SDdHX6PhTwE2M7y7PwVqvMq+JFXU82fycUFfhYo5djG1g21DEO9q9
VFNxEkBYBFonGLGXMkcRbrY9GvuNP86/ZTaZRgJAblcq2XYe0QtpzPYyK04bx4vIBBLH/NijjUx6
lasZygkBTkq8p+4iEJSsXICFGfusDFS4kUXOnC+a1UGCGgp4jbl+2f6EROfsrcQqSetkcgeJBPFa
6EzpZA7oowdB1Qqyuobc6kIzjop9mR6EgJLxFpcoMN70Ln0UelewFVrYT7MVTY8Kz2+yrvOlCY33
VY8/x9mQmSDCFqA4T+pEJ3PWfCOMJJKZ13y54ftbtfAG8hdIdzIVHvStvVYSF+9/ybnt05AzCwk7
LaYPMJxcc9Vwb9ZtqRFsWGWgDoeNHIt26suG70hANmn2/DKgG7YL19Jo44F96q3AXFpaBviOAWHy
+/GmegirRmyQpkZQuWvHxZZn2FqgruBnn9roiYDZO8SKmNefJcmTmxDnFIPDK/y1N+fs6bjyU4fg
3mVgrjmLAr7f0VNur4NzEUQSZ1OcP6vkMdmyPNNzW2ODABzPrxh21bnIGJWLwJowcnwN8ugPytLq
Ls7uL9bmnWJgRPIEWFshv4KB0H+dOA/y/Yi+rZOHbNpjqy24Ff9wLVjv2XV9DphRR8B6Z/DiFud6
ybD3xIQpH+KSBldK5V3PyK4qElioq4xy9NOc0JhESFDcmKWNk5QOG31FQG2VVHUvJ1tL/+KlBiqP
O+IuIq40iSkKgJaru0WhIH476k+TVBSCTqxAQV+IebRSbrMAmTP9JDSUQ2haQiuoEWNvxUn90g1n
QKrka8VJ7MBRbz+sXMlCWkaxODbQDQ8gbnbInSUGh9Tzgps/d2nz/WWO4tL3p4HuZIVyAGVuoasl
Qqlv5FqUVfG3w9F5tBsKK8xTz42Xm0hrLdYBA3q2gZwSpojyqdIRqKWCaNkAOyljnwFU39Voiyk/
VWwGNVjEDl6xpSGjteWbDhwGcPA+FzJMpp3RyXfkv0mTaQaDD/zR0jbeRrpuMnTpnq+Ias/et9xE
oDCt58DAJYnVD/k2H3H4FDcC0fBliZQT4ptFhVTu2Ef30APIm/kaUbo7KexXxBpprlmtFhdNDJKm
LtH9tftqWTvCdqUWTYEDe9lxphm1gr6qnSVaV8R9sF0G6a9YDfziDkpsyhzgg0zPMbiGwmLFHcnU
fmynJiXmvgw7oI0bta/5m5s5GvYXbRXNvyw133kZJG4J7e3S9j7XvRNN9fuZ0Oc0x8SjlI+anQiV
L+Fog/omj1Bbljo8yfbAsJ9XvQcS2LzRhRp0vPCNOLxosGDZy31IdzrGA3Gy+dxV3JrASt+T1yzc
/9xM4i6vOIqKJISV02z4XFSF7EVk63dA0XtnHdQsaW4hgemnV7Jyoao3NRUvq53JElLOyrMzHKuc
sLy/mnrORuS7/y2EGfcQ4nnXX4xP7ux6NsixMkWxPfFmAbOCpF1jzr17noaolpSIGloP//LB/84n
L46Yt4Gniyidu6aWuKJNX12e+4sPl8hF6m8yL3hLTtE40fr1YDbE/j4xrosqdYesqe4mt8vb71P4
GdnjYSC4HinaVi58cL5WTAsSOyC9cOr8Gulv2ByIGvGjNsw/s3pMKzgfd7tWFuOvfFs5IAQQQrWx
HKulA8oV4cNnYgHlYAh8YAyAxF2BHdYl9p5kZWffoEPlDl3MR7G9s3Lbk8WkzC4GSS3fiC1vzy9m
WYfCBlw0D9sECqWyc+1sglB/6CEDU+wv4VACSQ7iY6OOTc1zkzygRIqyIcl0p0KuDtThTKOr3Df8
Z/+4YGDbByrIbbKBZ6Ah/2QCpcNg6GT6ruPiNiYIROytYq2ZwTWxoVNYAdTeHBkItikjHTCKzzEL
UfWFcH9V3Kgio4W/qJPukQBsUTuVieo6+/aZ4GMEAok5SZMpY6/iqDBBx5scEMsRIFApBtPZRS+D
56JnGgMuK6kVUjxgpUX3tq0+Mihi4w7FlKtykJUgjVj1b4p8IdvxqihhJA8JZbNCmSFP4jaBIfKp
D3qE2V1nL1AWYSw/26cbEJqXZzOWOWF1ZFmQjHSaY5VwLG6QVMhsk07K8xaZmSLE/Ss7lfW1tN4/
5tXpF+fBXFLvH4dmOumLjo0arN8zROkHUIeFr56LjNs76xuXmgF72emF2z7OM0ZL0bTEpk38OD1k
I7tayFA2pmkZiJlZlbd+GoVJQsKP8GB/acFAR6/eV4xha+D7uYXfipA2uvfXBMyZLLrJdHXhJt07
IGW/UMfEVVPrLwb8NDvdl5HloN/oz/U25KbTFMLqpbRuYjp0t2zbPMcQ/reZ9k8sGKSbIig1Y9YM
ldc3RdKxVL5Yp4sz7+POUL8u3KKw6mcj74c7cTp32WgbR8vXt8sSMrqpTeG5CgL5e0xFvAa+6Kjg
v5J5jD3DvC3XMBbb08EyCyjCwqsLLylxEpgDHxSBXKtMldlmPxWFcDwLIHIWCE/JrqmT5eqnPxcD
/1giIyrllA5zAGERzRxKuqbLXAGvaCGfHJtiUZYBvBXXXUCZspflh7al4QO953co0dL5f39sEQ5b
hZSGpq/SH5A3hZTTbLgy5wLKsjrsRst9XDnxC1vg+tLR8Av8TLsUrNYfx+DmkDh/yoBHIRZJnfCn
0kb9AnBFE4Yg1CATIC/aE+TiTDiolaclZ1+AhhtLShSUDuqYVwyJGvJEVKkPOUIQVxfxsipq6WEz
efEWTA0OSRISofmjvatgQEQpAjBSOwCQMjU22qfL1imxwroUkkph4Sbiz/ZL7gkavsSuURk8QcnL
AX5pFwQwuE2F5Pvil+tXix78GphOpi0URFpKErdkqQtk/gw6lE1ee5/FAcf0DSheRkOGvOQVUlZw
IzGGGlRaUn4meaIy2bSQKUIB9XrSavoZe0OxHZCOJVWeXw5SxLZ7gygZBgbrx1nMph5JJzlFjh7t
5eZTBXJt3ngNvPORBwm9N44jlvl8cWGoeUdKMyZGANEEIp7A4iXJVY4TOPUWoIAceoHE2ZNadA3r
IKPzJpjvGVfogzrJoB+k7CapAj+pDYW6wKkgNjKjpjYIhZSpKl2PvUOAzm2DyyozfK5+aN7ievtA
vo5anHy4sm8zDRLYSwDJma+WbISa/EBJf8+UmhKmrUj4Ps3UtvTQV0ZJE4Xx6EPMubnL0pg/p10v
l3mTZrDzolmicC5JNERmWWYpGripdmI0Fo/43jBaKsd4o5VtYiNSjdeblutSvvIUOuCfZvdWtIDK
TsmetQTqd6KCuXHBbbxbKLbbGCNiPbJe/tMou8srY+37946lq/yL+Hj/kRJXP5GDhl4+07h1fRwV
Vr9PhDc07x16D11RXWZElNqFPfgvK+2O+deU25B9I5Er7NiBBhmKiyhD4Ev6MWnnbDX1D5Ih5UM1
+wONLa/ku9rNnEo2IHPhYSMMwASpA0k8CaIwmPl6W3NQeMqeh4O9t6Zfl49ZR85KP//ee2sbUvvW
I5X35mBo07YSFRdtuSQCyPfUPhaihUz5tSzGORPySzNquIIheII3uT/QiGzU33sWld1QBPJi4c6k
8KUbubsll8EKtNd3gBCPBS65cLX7V9OHirVvC9nPRR1XHgVfBGDC4ddBbTc5OPiESstEt5BfT72W
1hqIyXJNhqGE6rJqZwm+2QOPaHYSdI7Mq9ojvAGXJExrtebNcP3BWCpLe/RyRN2w8dY1L5oVCOOK
b61KzsQoD/+V9oBzdaWyUM+gjJFLWWKVsGugG3q/QavPu7xg2XxTXMz5nLBta4Mc3UcAxvucS6T7
Ft9mnUFlUEPlI3Sahq8ts81w4pRjbjHjyRox+n291DitgaJxmYcHq/zGSKwWo+HAbaSO1T6ivuKO
pX/9JsiQaD6nCv+RTHfPnMXoqTPrFgMY0OVOKLFPsof+eQlEBVOb2dogclWxqIR3nY+aIgyOGG8G
tSv+Tjc9Rvow9ikKzPfItx1JneBwah2BFeJf/hgy7rbPVvbhHHYF3vxF29Vy6GdwoYTODCE17RN6
vlEPc7hOlRBNzeB3VeWD2xjIEuPZ/8o5R49uheNHMXNPvZqxiQXnhrSyEzNqsEThf86Tn9WKPaMv
gcNcNJYg8e3TqQ2wYpj1z3sEeleOFuNkjTZIjn5pKX8Vk+bJ5DBgf3C3C9uJADDBeYa2+xtvSkfZ
S4GnoOGGr/BM5rv5s+L0Eodsp2scQVRlaERSpLqxTIF4gP5F9x/cKrdT+X6IfOz8UHnRT5hR4h1/
WePVuvpZvTZmsP2G+OUmXpDojWiadORBqzVvhNlfxAX8kU7qnkHAIHJRvRC6Obp7LyRaIW/e9K4P
1NpG3wetfWYj0laM+FGhVRumLQblu6thwCICCVKCrFiWQ1XkWoINMR3U86+f/Fmn9uu4LOxT2ynp
4MvKpPhiv2wNiAqc6ajnzjszBhDZZG6kmK5mUdxGNG68gawEZKq6chj6J8KCl3d0IjQtEuPBmVv+
8u2JXxErG8xzjQwuCjG7cWTf00/uTUTToxwb8PjMuTjuBzpG083R7hb+qfpg0p5EY017wn3gn0Do
y03VqVC1MOGaQt+v9EVwV0OEZlK5AS/V3DxGKTLu9a7WudjDwDxuanRwHXGJiy2N7U570UJJKzSP
X1nMZzVnKaDvxFdd0XF0KYQIZlEGIRTHl/YKXXP/nwS9ADxhjwKZ5bXTIYzidZRRQo99e6XzlhNM
CFZOdTovnIZmHZsY/FwMqJpGZ2E0LPqvxtmQVlGgjSNvV4zfnR0jSV6HGyZ9uVREQXbaldh0aoCV
A6J5jcWEOQBEPPqgQmzDu5xQM7o5kjlW0Ew4IcTahNz3Wv5IOoXu0sgJqfLHjtYfkquVH4ue6jC1
VqA0qM0Eu14Y4Z+kkL8cTVkXwHzp5y7HRGkIhkwTesyjwE/1J0XyLeDxv3XMSIVRklpufIuhx+RS
H0CSQmLPcu4YrL6Vwm8SLc/SYsxG4DttBY++4dlHNQJrguP34hNgBHuSEKPe7opICthckeRlKEj8
/xI3SkzIM0kE9P9DqJSSKKdDdWeGuDmKEjF3+FMIUCMzPMvbe808xa56mC+yEwcLm4TczZn1RzUZ
TEIB7iPEIt1xFGB0P3PBZDE23ga20uTejLuHr/COdsIm+tCEaQr1kfBBUrkjZiruQU/MZw9sFF4O
JKXszlK69mVktD3Y6MNQGAoNp1EaFthGr13WCT4hA4dEeF7P7az3nDSXhQSPS6zTAvUZL1q8kugZ
3JsUUl+B/H0zRNkt7lh360j21H3K2b9SkxADWvITh0JCZOmYru5sQXw9fZhFdZLrNBD7uxdTkbvi
/7ADomiQa/Z6TYXvOStUwIQOIBBXs1iGM2A+egNptsYSt3XgYSnHPPyb0Y5Avsy3huUGLF4Yiu2h
tn6+gy8jrELV/akRID7UdN5q1rgW8dMQWZSkkes/zL6F7iJ5KELQ3t0l42F/y5WPyfHS6XKKJLOn
bOaUMNxv1NYZqwxBZ9aPdt83iwp0jOoQL9WP7wvQWTqbPGjKsYpkPRZk0O0WX68ExfALy/n+EQTD
7HOAKps87SYtqIxya1X4KOwfkv1i33ZhcQuEPdjmJwKglY/YFMLn9gAowSm3Wju8tKgctMljx4jq
BsMxhbkW7lPeVHz2PK/jnNKbvsOyUXov045Enb3Ip3zSPmZ5MCfqSo+eAgu9k4PAFIYD0iCPq673
00Ny8Ke0VcrXkcmt+WHPBYvTjcGgZrZqEQhf4Y0vxvxo9gu20LAXlu9I97Q8RaIgEDw9/eH0dkxl
1uDm5G+xmiJ3KDpq/cjoqPcQf6DSY9J6HXDyKKd57Jx6B/wjRDDpi0GYayzNn8QBkAAiKDXqQCV1
fbwKfCO1lZhNqqoUuhoV3aKMcM06KV/rFLy/idWD94Qw5E2rGEC6eJfiZgz7CNmNiVhWesS0aH9F
s4eaSxLpd+ZSYWonk6JcJftb9V7xYAMBKwzd1PyfKK7pRUTi+fhh9+QwbfTFAa0HL9TA0mho9KBO
qzeteManbNyz0R59BHgls7TvsO0rxsxNNM+aE/BFFOMUvwlUQF3Cx1c/mH6QKe0h5R2iFMHctc3X
vytWLfzOu3fGKBZZIT6sM+vm4U7kSk7CbsQg7cXRoC8Y/7NjXmOOzZjg8d1WV54g5F21ea8lTohr
s0byTFJz3dswXT+S5w/d0iYRBdJYjWiah5VCMNgTbH6krw1fCN4VT1CBTQNrv9sosQyCl0vECAir
wrl33xSuP6wHSWQRCoXG9wh78UYDv/U9+5j42rNG0bKductr5rFmtbDB8WVjFSSfQ85ba3Qe6pSR
r7/IZWrbDlSaHQRGmy1GyFAptfWYYVp2hxKSjtSsFHxeTPc4GkVeZOg2RXCcl+yvwgcA7JiW5zvZ
Q9/D1QpcJWWuBS8UqKQz0TzQAAAfPH6pM/kxe0C9oBtqI/oPHRYZ8fAchqiCt8EWw5H9qu8g/T7u
lYilmHoIO6054nFG1fc5OHHfo1HeCHiNFMz/XSWcUb3MIvQKgEyq2z++0nNihjbk0aX18Ny+PdfI
sTQZRcXAL8mSsmyH6c8/2REDKsoWnbc2mAuwjVIjLpK2oRR9Lj6dUpybFAfaaEqJZpNcbxiaSoXc
OhJo+YkM4FM1z6kkI5LSCs+f3z3EcjYbuJF8690TNl/ErMgEtSPcldH56douhaclmpX+yjZo+WjM
K/Cu1uCBubkr8JWSvmPZSnU40wA8A9vwTiNbTNJFfjxjBXqaqbMVHQt787cLhvSe6+ZeZLzouIP7
bQgEMccg7K3W6BkrS/CZgZra0cIB9ZEtyEhndf8PfzD/xSodKTd1oKqJei1hiyUplZSlO4guyLle
VFXzknAgB8U1CkYd5JHZG8jJogh2qu/bAQCsUakF9A2t5cLocfMWi9xPcCWsSECWXhBmiHB+K4PA
+G2pn1avJB/mYulJ1mmNSXmVx+I+1x9g6ilGri1myNNdGcBkOfvSJQ6B9zg+nd9IoT5siPPW6Fug
+nWhqe6M2tQDhlo7QZwPSf+8E9ogXM9ouL4FcsIzDXzCyc1dHK40uMV5Xz1cx45Uy6x+XNRdZZsU
z35ZsQe2K8DkPeYUzJyozPrUUCG4Dk/G5pMXCbFfPt1icKxWb541QJfnP50t07VXHaycmZHqLKqA
YAEbkPcohYCgq0o6OIuNHCKKkENhWQ2MJxo2Veh4EBdtgcM6NhTm+R6dcLR/gcAmEoJQWR5GnvH5
+fGttmbb6LdI+zoB/oMJX6TXm6blhnKg7qAG501sfYcvve+Tribnv+AJY4kqAFP4+uvIm9Qmrx2/
adPBqqwJitj7hn8gcy7yCJNi8HxUS5gWS8x9FYdo81YgDuLTwrv66fUqYEvk/v3IiT0kD+9yNTb4
G2dfgAdsqeRtzjwDWNFrPmqdNtPmGap60CaQ7ktX+zCvcycltkyLIzwhfiTC08MNtFdaOYny6u9z
DXCEA79AreWTP/DTl95QAw0Yz7yURrK1OCWyM/wnDDoSPzEaqWlmEgTbgQeX/e+A/QK14V6JnBTL
dEfPRBl3TohIDUF9l9mceNlUNWKq/E8elf5uvVDGoWy2Sd8UK025I8MOvK+0L3ndTjRBNhq/u8Lc
fv1IqeHmGSbUUnSdkY8ZL3JiNyR41glY+0owNHKEp/YgN7lcGC7gPyj/LegdFnJ0MIiAHtUr4JNb
glk/zZKeBYIfJJ2MktNUFityKxL7O5X/1/17Y25Xm8VlyoC6uVfAvsxFBES9DKs3BNLRvBKJRDlc
aagVS7U8OAAIJE96Y1Kh649Xde1LH0gQKhwKjCZ9QIg8HV4MkKYsauh/9CfJS5XFV0t3R4bYFtCX
TZya6bxEqNE6v0gj5hlRXNDtesyzXPzhpoJGzL4U9ZCD/+pk5SP9w2YjV5O+5zesaJM6Th1lOgTm
9KmrEJptc3efborg/8r31WMoBHROo4ArYNKazOgOr8FBMDtWFRX6DK/keP5tI3diFIkRAhtBBsQh
9E3WFTJ5aQq1Y6PmtpG7G0mupZtOSIYR9IWsB96z51jwC5eN+zi3P9zKildYC36i2WgLPEH5oECi
yCdWzK0pOZdovRJXcmJYb9bakF5Va7xwbfDgqRfk73rGLBRFvN/AjV5hlHlPfxPaGydrPFbeVMiC
gDI9dwlFyBGyFgkHahKxWZFYR7VzCA9Q5FfiYi/Ir5hVCCdlB16Wqs8tTu8/93NFtmShW7sY5jlC
CmJt6U1LpKX1+t5uDQFszTJHIcVFD5Kxs0XzAaJtwIqWRlp0HCGZWUnqE5lMobfwO1Swl3wmfIyV
EQCv1O1EHuYXaiLEFKsqfNDXW7tJFuqnb0ijvL+GHoPr2lg/oksrH/DYgWyedRjTxlJVxWN/u72a
IHNXi06WMyGROiJ/qpBw53u2j51TOrx4YmnfwYMlhSE4tGl08MdPxN6XTqXHwGfUig8+NH78jfoh
WbbsYZ9NKJbDSdLaWXJwU1za7/Ih9eODWA3aDSGTQ2HhL+fZt2yrMk5P69q7nwMz794TVy6TQu+Y
eaDMEEsToDof1g5U1LOxgZNEvKc5JCst/kBMns2agfjrkH7STtuhpAgx8dSJOUHeoSiWCDdIj1+9
MHer8CHZDugs4CUEPg6+oh1DMBs3Z2kp04sS3lRegkH1cFDxSnIV5va/5dBFumPbEZ7vgsAZ933V
d5wdboKmsp7LN4PepQwmiU66pzgDB9IK2QXrWaBz3+dWxpLlnc2DbJI/izZk5TDaKx3cyTgHgsv+
wPTCgCwftZIsaVaX7fUFCEyWUehpJJEBOKazUeWfiomRcEdqQZSZAN/yV3nGY0Ry3rGpdDJjm8WS
mT7Jw8rl5o/IZMLuvev3pQE2xs5EZuBW3VCOfBsb4dQKPgchVS79vNbMzRD3rwI6F7Kr1/ok0wYf
1yvB721MhGhJ0voX/j8Uorf37IBCTjufSxx1AvNwxAqqTO8ySUx+Ih5jKAJhZuZTyO3iwevZ7yf+
E93p2Kob5YOW3rtvmLgdhuZWD2dC8kvPlkTz4c9o8xziN82sDwxdW4pH7dRC4umKV4I8o+Fnt8sV
iwdbG/mjk2UjFET6K/gyxrAzmDGB1h2YHRIIk2Hc2DvumYW9M/5kUR8nmbL5PqYhcAavf7tqUzGp
W6TFAPDRB3f9Itd1Nx43lZyfLShgCwWkePEQ6WH1RmLnlRdAE1GCj3IpALCjVZ3C65+ksFYUuY2Y
/DoO4rr32KSnEHE9Pg/RxqSKUu64i94fg1Xo1Ww5cubXfxP67pHBMCgDD9Vul/nxYO4ho8ZKBc83
Qr6+URLosEPJrAG7w2++F9W8JEHhq1Cu94fSbfkQ66EWJV+PUfpHUMa7ZYLOEtpH4HHwd5SLWtAS
/JMSBPOlPrQphC7Ysf9AXKi6spumS3MWZULJ3qNuJMnK131O9baN8ZC6+xfJ5cTVmHYXBLUouJcI
r/3H9jl+DtH+inhOX5vRRyy0IdKV7cRDqPqAHBbbXHqS2SDOXU0v9Cb0BGpLdk5njagQWJy8BE1u
1ab/0/0y4rr7As9K9wiC+Is+7kabl866VuAXhxkttpnQ1pPrR1O66CIZBftns+6yrFyOgGJHXdNr
z/W6yJR1JmfpZcPWKYm0/sIgwLP6Ib4tUk22bCCtPGdPZwdY3S71YYjv92u4iCP9NjUzqYhNI5lw
wWqabeFdWFfjABfTSXoF3Fis/RyNMVO4ZtdEPS8gw9wdJ3NVQs7I3xMNQ/XCE7SwpdZVh2+Exh7Z
DhT/+KxXsW37zrtqpu0zqY7pW9o2Q41bkiKo/mR+I+0coXVuiOW2hUJ8BXdZXH0W/rHoNEAVo6y/
ZTbU3GV7yzurOGrruGyzWKDVHiMT2H8359WEi/XdLh6c/x+n46ZcPGp9SaMGjPKlZtmx3Dcu9Pw0
vNBlkF9htY/jflqV3QKhA0aZ0K4IXu+OcpBIMgR7c3IsZv0959vPopfvqEzQI/YqW5lm2NMTj02L
WSYA21OxMyYWuWUu+5kH/uQIdcyWza+NBbHiG2a5//jgePpZnCZm5uutn6OcmoV149WPO47izBCZ
bFzNxVBtvS0/Rgpt5dU8H/ppBxJv5PMQREr6fvb6t2iiyK49jLPhP6EcJdknWjwpXWmoWsZr6o+x
CCbYpq4QVBwi9anJvoPGPM1+aRxmP5IgZ17ooVAPQ/zzdOuhuLZm3X9db6dG3Wq5OeeJi4ABqky2
w2njBB3B0phbyvSgRq9sQ4ghQUoelMOaysas73O87CQJ7s9HRStmyB6Cr3H4Ws4hQpDwH7JqjJeN
kzCHpDgSQQt7dRSk3fXQK8uMLg3H3z2WNKkRoFJxEwacd78mZhlWqb5XZQbRX8+7Flal2luGD21z
CvCfVdGi1MpcFaBriNKv0OcWz0bDz9Q0fCyVPf9Vo77AqmXMEA6DuKcwOgWbPmTrW8h5TKupYGTQ
EqD12WmOie2UhBjQuDpgnrMRw+5PrlA4MzFUyY63pRXruUfhpjVEJN7FO+3dPPT2k64HGRJVxUml
RVdb/BAXIWo3JF3ELpCHLlLGlPV5O8IMh8v8A8dSeEI9Xcg31B4rv/G/5yiDStq0V2TcJZ6G2d81
ib1mjxM632vi8UZhU96PjHn8cJTscIKAkrH/ceh7yEQ+TLhuGv0t+4PDZDNf1KH5AnbmoMk0/hq9
RvBlcKCRjC+5LGCO0uCVtAkE9rRttepKacrewzHkyOBNRBrfzVn0N7xFaoRI2IWkAhRHiBBBTrq2
PRX7Bo4KJrFWeJ9aqi4j0zl1JwO00Kkr0TXw+po8wYeuOP6U5t3WSbID7yfrr6AoiQUOeLlywxuq
hAm2207VtCoRET1sky4QW5xeBSPBZVVzUpzLl1z6cbUwyuxLd3jW1xtIBMu85SsqVRxuzrkOE0mE
qt7sN+Or/nvTdk0STGeHmyvBNBIUogGFYLT88YWYsUGO19rjf2mNfvRr86l9wxq1Y07ZcCBdDt3C
fJhrgOPAr776qHxnmQFRKvpLMmb8Ypzqay+XDEEr3z8iRcYSMlelHisVoqorFlP4ipXNFwjasTy9
zgwbJXLTV6t8khs8wsX4lm/vX9B1YUhNHGepr6BOXhg93E3OrEaFVZA93xFnvA0uCGLOtEB7DNXK
+U7grcF7MkMBtXykyhnF2fYCm2bl3OmRG2YVRQG2wfxx6rKro+HDlksSLCA0ObyJnYoNopz0WfsR
bnhz47B8OpzLYVo0cTqYGPAVagA1ZSGXKttg97+vDAZBXDj1Eduf7/v4XdB8+pBtoCK5VlWJ/8uW
i31rgyanQWHVz+cQmEnLg8xx52mn6mYa7ieMZ8KmB4JzL8igkOg9CcV4UjSbb8NG5a/o0hIpZui3
oUX8F/sz6VH+fayMnPPSHCiqPoGD4+xTrvN13jIJnr+rxn13wTMlUitzfF8z4E0eVkxO+9LOk8b7
uTnkLf0/kkhLmn3iv5p0WPFAtfumyYEAXhuALWQjLvFx+zrN1hmEYgNlU0B69izcKznvLg3eiK6y
rNHJ0jrMjicYYeD846TrlvixTv+hnLRxgaccmukB1EPLua241haIzfB/JxHLmuToSy0QQIwwOEjC
GOYxxNYL9VDxd9ioEkV76fBczkapvewMIAWgQSP21uDFTtqjiokbfKpMjFf7Rk1BiTEHEOCEtBx4
NPwVANysdajGKeAA8fuoVUgMK9aHg8QxZxAyDHA/9oT5rOwCSVpIAFCR8tc79pqjIakuYT46uzH4
7oDiBzvRJ/rRMRZgKF0itilmxnxi5ydKkw3q7DpJxaY3iCNr/KwUUNYHPnNVQR+WDM9L8fnDN1NS
Tn18P5uG0b7lBlfbU3Uu6w2SOAwCKUIkF+h2vDFEEhuq2vDn0Z3Oqse5RlHj6uGcibr4BAHm1wVJ
SCntEYrtOVWmIivQJvMLnmvpiyuCG2OYG7vPE31rVI4wsiXfxWqVFYWvArytFL1ACgwbnSJWShbd
4I6GIu44YHPBAC5FdPFVCE5EcQCCoiVZBZUfEzblHNrXAS4hb3jRH81B0U4dtdqeKu/VcVPA3tOM
jfnM1JJfqdOYffy8dqbwExWRwwYoAf7XHoW7DthNlo/HqNRsH41ZB19+HJxTRr5RfPJT0EJ8apb4
yFhTVty8MEoqhp2WwwfKlhLQJ3AHPPVsYgPpxgcrue1iORxAlkDZYje1WRY13oTgMxm/PDCJ87K5
E/7HyAFCzyZ1jJmTpB55JrktOaHvOm1t8s6r1ALpjy81MZ3eTGdN1aKlWIbx6pCqjKEig/BF76sm
d191tv5occVrMLq3iuY2BBLiMbjewDQDyv87g21wvca55QrSL0iix3iAy0sRyzugEpJSjUAYM8bY
94MgQCJeWj+xde+b0ydWw5NqAync586VibmbqMby37zXeJBHkBuiQje7cZe3/bYDr6gSpyfM6rXy
OkKSTJlO+g+eSEji2r012wjoJNk5fLWEC4oEM0UEQp951ppBtNRGktAjPTZ0vnx/6ujIKqf0w3os
Ms/J9kQW6iEIyqJC32YJg9tt3kH90HS6/g5+ovt2R6oOefbM/zpwUjqz3Djr9nbJrSAcCF9QUSN0
CQtoXAy1h96l7guslFB2HPWhUWzmIWC3r9wwmL6pE6jps85Bx1yu6IJ2YpFOKw9uneb8MtHVkVkc
UXZVUsrFfpl174mKCxpilvZLIaEiue/AFGgqcDRQylHw6Ilpwj7/y7ltE4Pr2/dTRqKWVkzKN9v2
F8NEQfdcjlBonOCAYOs5wsvJxqkL4reog846TOxZbog+iarMDwm6iYJwaU2NiYObXu+7lXylgJXZ
HcahcfjMFzEwngA+2TcE42QoL3yB9qmCuovhDw5n5XVee6KYBoT8xP11TlkEbILf4aGZUh3Da1Av
5WBwXOemjnJ2m21cO8lpCBVEH1+8/Qi9GrgHum5jXj0UZjtbQEsVDKWXlFFnxwH/6WxTKb5Xvn21
SCnisbUTItq8gBDhOPVPIeY2PDfQeo44VrXVChR5X3c1RnzKxF8D9DuegblpFOWkeaxI3EQ463FD
MgmXn+GpxCbyLuOOkw6sBM6/QD+KZ4LctJ1sQ/YcrSLsNXsiuOAX/ZcKbMJ6wTvk8RJRIEqH5uXM
gVdo5yJTMFkUj2wLNVKmbsmJCzjX/XrmnGayFDQj0X7skMsBAa3pvjVN+n1SFn4B16RLERDzjzrd
gTFcXIyO+Kap74wIyD44oPLwl0cGwqdC3LD0ZSfJMgRaYFYnHccyrkPgD0nWBEe1/iz/6YVXj1Wk
5h9LoVvp5IzH9DtclYU8uvxqd0kKnHIhT+4Btd4DancGGKF3JkfXZjqhOx2pm2m+bmMB3ah37ozE
AMKlb6KB6A6YYZz5IfNPTyhtQiuLcEO+AUH3FysEDhImWZ+p2xCnZuMI91Z5gNv1a55c6WdaZbaZ
eucEgCeYVRvJtQvblnpgcQXw3y6T6GJ5zkF7j6wjBRIPeTHZ6G+oES147hoqP9VxwUgUY1JlAy/6
JUmoADbwKRTd5Owz3b/4cJUIxc4y8wVY8MRa0ekXP9sQSonHxClG4LCKrlRYfo8aJMikN8t56yjQ
QROXVGmDwL4z9H7OQghHRb1kv+cwfqGnmNTkE/wBqz9IFxRfZLjmcAGjx0DU1chMmxpiGYmBOXcM
O+MMkmFIxpSmRM9ikXjz575a35s6Ya1iPzfmyqL3aB2Y/3JG7zrk6ElRsJZsVMYQDOe3kqAojxEX
0nBKGKFmJkV8c0lhkPlZwSB4cs1juNvzmQXp0MVp/+sd6OgL1XJ2GpmNS50n3bXvoq7zkoXJf2sw
1lhrY7RjfldPYYFYbzvVTZDT4NIb9anaWivzhQAuPYvWvNltz7+9rZ9XCEjoMt9x8wkdMGq3dFn2
t3ViyWq+j9dIV00zfFScdSB+9b7LiW4WHkLqhyXmdYyPMnKzxPoJOr5YsoRpBOnFqfiilmOeKhHc
yxQWNSKNI6W2hcx7i7z/awkuj6DW+/ulFfcAey94mC7idaojlr1WKB1gUcd0Zg+YwpkX+HhEa6k7
bljHsYhLauEHPi9ASPumkqaBxzJ5iPLD7dAD7+jqXSw7zGp/MQ0LZ0sFFqeWRPvPn+gMi5ybHBri
UAkO0zMjrrw8X6hM9Cqy9wcZRQO9Nu96hHlQBPA5gy27j7i4aZ1CIzMsmVhiuGBf+W/ucsEx+Gv7
cZtwXYzo726xrPW5h7i/XsCHH1BzgMqaHwpTYVBi8KZcVqrygJoDcNFha+Vwtw+1g06kiNB6aWzG
wgkr6tQPaOMmly2+Oc0rdFcQwKA8Q9v73QCWo2UHH3bfrNeFR2K5cDhvEMZRF1qVaHdPfUBjm+Rl
H0UO3BABxsaDuA/cqVIh27pUZxExaCD4bgt31U2cgEEUl/5rMaHnPMnAe/4WK/6PXRA87ddcbWxQ
9bcbvlZb/lJ2qdnI2K2B5lrGopBD0lC1vOlNBlhzuc8TAOs3ptJ8cIdNiMyGV3yeFw6IdhiLO+cw
ScSWwABd32W29qtodkS6QeO8RLOZvVXCRMLZgax9VlIzp7k/2OqNrWMNdlvZVhHcoz6/zy6n+Fe6
kTUBftFW4DzJvXyFMOJKlzFJ8KNyanvbyh8VqxfztuijWd8tMSq4L4wg18jHQVI4mNSsjvmctjPG
k2Kt3XbUiaagHyzDpymA7D1v6AkystiPHViNFQTo2mG3749XT5HPqzLKPk4VBUsbWHOQzYTSmW47
XuBVF0KXO2vvQrynClX2kiSWGYeOUodswEhzuZwnfNumyftT+bj5gb4VzjJI4k7q3qVO0wQmv83r
tw3x891m3aCPymcdCcpbiVpeGYnY4AXT/kV64XpQvKJqtheYA0in2mJkOaYiSnAOY+kjPZW28sGK
UfL6Y5xnOzernchxxtUeaC6CybkXGflfeOcnKTgHhED2B33mIGItrlNLd7zVk0rTjTGXGgrJjpRZ
m6rPfezF9KDbSSdK4KvVC+Sa22PHnj3Hr5kMOWRbqaP+Mx4dJYDUkLdyBwqrTVNfkqcNMmWbaPI3
T3ZpAYBisFW/TWJOw+19TMGgD0GeX9c13L5kJElpXPGWTF07D/kPLFWigWR1ybcy5qemyhxMa6rv
ewyptTkKB11zmy03ZC9RQD+YYv4QsrW+DYCg7MYK6XDXXszSQZ2tWVVvlIGI3cNQus6e6LcbOj1u
27zgeBzRXJD9efX9r2h1c3T8zkqEylfXhPXgGCsogLyikQyytR94HqNaMYNSO+q1CS7CmOXwr+Rt
keM0uWvgK5hGJUeXKOcbVtesOJOM5i3T9FJq+ZslAqjZN2rPXbVVOm/sA/u/GH5fPM4X8ZyVrpXM
Hxa9dPHj9U1pL5nZU3gq/2aDz65sqcuWIhi6i/u+BJqTLvIZqzYuZXfc+LjXjyWGaVLRcdV5BoOO
SBZojUDS0cJdoUiHqniildWjTyooW7CG37Mee/jYW5XicXOT08LZjns63voD8GcqSOJmZox/OXVL
kHoGtlCBRmmMaId062JykE257kxC4RHQkkR7EZt6M4mqmSwSLcRS96/eyLQWccL7VEN824q4jSJS
YdTbkKb2rb9IISH1OL0toUlZFKUiZilm59dXqoBeKESkab184474736O5c1H9UHsj/NDLLGuqqPx
3scQPeCAzVIpo5pwJVYnFCTEV3xvZor22irsKDbI4Ty1PTVpvLq5+XqUF3ZcU2RRk99w7L/Q6j73
I7BJ47lWcQSDvFw3IeOxY+VC2snZ/3zpmPzawdjrBlbAb7g4FTMy5TBd3mTyl4QcYh56k+p8GO42
/IKBywCfQ2fC8rz8hUBqxjs5PCIOhcjqnIXD3g3pNnDddfeQ7bRFphKPIS2i4nYQ5fqNJte+7iXS
+XSvA9tYhGqPLizxDt1coZ5jWYBi4KRWv5cnHXopqWf+Q1tyi9s1WSDv9wpP9H0OQrBlQ/JhQdTM
O6l5y5vMA9pPdiACxvNc5sfXGSby/eUwieJPa8FJEEBqxptuQVAByZhcrpRc/PF/eWbMZiZI3bwD
GYmfpy8Y8qxXlwairXKuNfKCWRfSxqUf1yYvYL2AgKzFoNrtjPR56uD8LWwn7t+12goJU6RaBM2t
SAAMcNdlxluyiy7Q9VCU3yps19WTWzfySgxhTkBFruaMr704ryyyZsO63T5jfGaHX1ecVjctviWF
0pIXMkWDx6q6PxF022XAPtpzt6Ygzjx1kkaafl7PPouxhr2vejOTcgVj1NDv5271AfiC9HnGgcer
TJPw6YpaG/9jO5wlSKG6/bdqSc83z7pXepXcWZY3/f5YNVfKeWyGda9hjbapUy2DqxnJ5+rdJ8pu
zrUI8fjQ6hPJyQkwD/oTV3Oz1EGg7Ej0BG3E7KnrXZQQuyTHyDQG/sfdMtzxizpfPs29tL1q9G7T
ILyskhoRhVjtfWllHYfMxMpMIeyQha776KsU9RqyJDQXsTpGJfrX6NoZiwQQlnuvjawS8CnpXhqR
kNtTWf9NTYQMGCGXW3wJbKjC9o/pRlhtzFyzhPVxsxmsq96T+Ls80Sn+0TCRkWU7cmwWIevfm1ov
0Hj2jHCY/09rO9xhCXSE1K2xmnIMFrcsPp6GMVNYBBswSRo1H3AJGVVjp725MqIVf/idhZEZanFs
/WaVIj9y52Uvxcb70EsbcL7YuDi4BBDgOtq0HknAXlOA2k1JO3ngmyqde0NL7RZgVR/0DMYOm/vq
vLfDSsqRPAoFfQEcxawYLKCj66RmlKVQrzRZMx9StIEEWMNOWoyu+0o+mizg/5r0Xw7INumW3BzT
ZHGQQ4jbKWXgP6AAunC81Hk1vQHnwc2LLz730pfapVppZ7ap29525IlZfMmO0jhfWmYvxxtuLMxb
9B5A1m7/vz6aaErJdQ7SjcKw09exTmQUdRUbIKzyuGWPJYKGSeKeYWkJvNOTzhdLF4B5/KxJA+wf
jAWIuma2/Ki7WSrkipgOZAs6UNAnNLaLuGoN3LP7wr9QEAK7ZfpzhQjCWN65qQiDSfMbW5i6Iczc
aVXct1Y4qQLNvXDo84VSDYpqDp67TGnhio93tzTBzXKNJ2tbAGfAVjeQ04sGgGtYf6zhpTL3jDFX
mAT9uUivxQECxJmO3cSOafLEuDi6slIbBDGf0XGD6XYrjWigMykqB9PKKt66rRCIQAovSYUfoQGv
ASZIEvoj9GYMQFHfHp5EQPaiVp0LnE7Kem8JjI584yF5u7qQHwuCBreYZXW8Gk1ENWM/Uwb2YKid
nJiZ9XsLqT1v4K00hkBHMNog4V8TsliHjehAPYQw091A2nBcV29+7k52fJz8dmYPR2jvG/phZvc7
0s1+0Oz5jMp27t0tQwseONDVX6m+QVyic4v7f2kUZkvrkIj5iz8YLdVJ8HxLp60bNNJeHl7CTWeg
v7P/xIZ1P4kp5IZDDVSDxxaU8MxTlouudoum8PPVsefLlWVhceVTegTTI1uTgf5EsjNPGGEpEDy+
r7Se650Q9CT1dmJngZI06e+BDZivxZT25p2QiwuR1G8n5N5qOhjS2aO7ZKRF3AqWI0Lklai9srJD
7QepNasAraNWblGfyPRy1+zPlu5h6WeW1fvnHNq8eVN7uHHI45Ga2COSpAeTWxFj2J0Y+du3PgrW
G0f3sCTAmVMmTsZSZDqF4jRNUIa/8LMBFtnKJEgjF3jWZz+ZY/FfgK9AYuK/Tl4KOAkxlRZBBxQd
mbj7CZ6S6FaN1feYXumf1Vu4alSPRefphfjZXyoG14lYqUrYT1BVnf9exAnYV24lpAD4VqM03cTM
5JJL1ImMWcqXiRG0u11aewQnajUiVtze6HLofVzbmxBhXOH+/PZf2W24o5HMqcYHEbluuC44VsEc
v/G4MpsLi6IDUzh60/T/kor5lJnTQbdOU1DL2nmaAxHcoltKM4FaAmN5rH2HthnArbwU6Jlk7fo4
D+/80Yhwl74D6AlIYN6SWp39/lRJKLuDJC7SaQjqyuflOuavkNnIsVPNr2st6w+5IoZlrCz5zeqx
qQCqzJwc2USt2d7BmkhpyMLeXXkBTBVwzzmvyr1BLychRK7A6ig3zu5Xuepk3alvo7sZjIha79WP
YKREyMkkaEcnP9YvbONdcRy/lD4Io2EnYC+vSMkh0sEyp15RovSNJ9tQ/VYGnXjrtVENaO8BnBjC
RhW/Ep4SDQLnnQVmYkgvPMYyBCCJorb54FraOOKN+jSNnYdQqpi34yoagblCy7orD0OD1qQJU+hJ
j/5sNhkos6pU0IAIV3joneoUaT3HZABVMufA044TpS7kmc8fTl2v6yOFkCFSHWGL64KtYmCxwBP1
sofL3TUd4EufoUfWwpiTQonuUCX9PZRrxN5A+b3Fo5+JYl1gDuPpXxsd/+OhGIwfQDaF1yPI8c+v
Yb3t8KaY90v6Ly0g7MofDLsBeqLNBlpIELXPV5sA6UCQvMAIz/ckfdRY/KkO6L2/AVufVSDaVu7b
lLc8zMKbHT3KXIoepdAM5O/V4ukU9FXnNZDBb0ONYClUHWXjYHqfI3+n+RpzkEeeLN1oDunxf4d8
ew+MvMW4aC/fW8LQ8S/YdmO+rL029ZDIfLuAaKGCvJaZzaO6z7uwcExY7sgghvA5+GKZhe4+T8JH
ReM3zeaacRt/wKnT1cCq62nxSTrKZ+yxlLkTQmajjK++Hc+kg1Q9B2M3OdX8ilbRLXfHENng8z7G
B4luTjudzzU5cBDhwHNDObU6qH1BL5cTmNTCCCaqeLkZpcWNbvw6MPerd67JLEcpifNQtT9D5dWE
cyDIUx9VY3CphNvKzJdMXrAdYI/RZ2rV2iKPZZohLdXdZrCBG0tdaEZ7M+1+u3VqUNwYL80ydeyX
Rf0Q2CqM2naQfBTCVBFewmmCKaENcU1yFI8YeOw2cVo666C5DGgxO9hQjdEKTIDDF37EWsoMf1SU
7ghnWovuEBjikZYBPO2MzaycW42r5Ag8iXmj5knpdK480l15+SvSslGdtn1tLGPn5Offu0L3qd6b
DlNaKoH/4WjOBMgQhhJAxcgKoOIjgefqijocg+KFrCZ8XJDKSlSL3OhprxM23lNyv2FPIc+pd7yW
OYa8k7LaZwo0VuWpq0ZqMDMj1Is83JAldDidBt7YdePMDis68ZydYugt92Wt3yfqYRZN7ixRiYmQ
YBM90gn1jOWbllCVWMgm4g8DHEA6xf1njf8zntn8Yt03R0Sa3L7M01GSDCxakD5g8tAF2y8iALdV
wkKy0ZIaMFlGyqSyOfWuhZNcP78cR7Rim4Pwhf33O65I9e4d8bKnpNe88KpEyi9KbRUwtHEG7dWZ
ZGQiKtkXY+HllnDxLIFdfMFn/XcqXjNQ7eNGmblRTd1wT9qTERMJAWu7NzJ5yaitBJpqvnbtWg4W
Od8KYd/WztgNoZ5hFeBRVbAYVUBx7MqlF+CHqWK8+CAmZ2Z7wVQ37/G/U/T/9XcY8jS+I95HiY3n
7r0pn4PDQSAOO7O0bQooGEYAmG4HtlO0a5aXjgEvkr9VepamXrGWL3TqPVn7NL8A8/Yx7zRbkkQ/
QLycF2nvS4tbUs4n1r+pyWCBTiKxyiX0ZQ2+1P7tIYSyuKdh/+v3wage8TYC8D6D2DFx1N7EPIOI
XNqx/ssW37uZeR++OFDDnZ0KGi3pn4gj+f43l//WhgqcDB8mC5wF6loOS9K7LUDe+QIrsFj4oX4c
q3D3eoECSE3Rkl6hRHF73GJTcppVi/uPqOkKl/tNwtGs6vPxmwb9Gh1yS/TenymN+ZBb0ut+yoM5
W94NDUDHTOF3Se9/9VuYIt/lyO4SpEi02EBP2uBrha9OLC3p9My5jbJxCL+hVyEXRtP2kat6ymOg
DGX8P2VPBHy71Nr3tEqKwBFY2gXQF+qxCl7syQv+5yfQP3ydlQni7IiJUukVKf1fONRcKrZJ6aaP
oH1WyX8Ad1G1cj+Z9FBahNR/sjb9C9UJrcTvfi4yaQZx4jAtHJKmHj75OsG099Om9VhwPiImYVsS
tLSsjkOcDmUDj6ObcPWO2a9BLfP5ZoVI/STXmjh6xduAkpAxfCNpH57uQFzAlLjqg8DLBkaLl/Zw
EEAzwf3tHlv4tyihRn8Dzo8DQRLPYj8Ic8DD+pscic+4SCcEh2h+4qXsbCznuTGtukFYpfvo37o9
jj1Hhlab/0YSCYjwaax3f/a+2n1//T23a6eh4ylKv6DXX3BGn9iEACcoE1nfL+ti17zoSL8wUSj+
alb8SNiELgKkB0QQZg0lVJ9ZZRQk0EYd2UyR56PVKJ2ryw+lE0aVQvk32PwHYdPfzBCG5R7pu2ML
3Rp78B3iQSRKbjt/WgCmn6sCCd2CXDOyVW1OVgqIhuzl4Ddh24iTmE5G5DaA+Zuy1art6oP03/6l
Jp3RNgFtC4t/T1Ck78u6+o7ANI2jAX1yp7HhxMBCOKQWuCIOXyEV44jh59e6uBHPozg3mIWEP5r/
NHFHylNb1qz4J818F6LYxCAmDEEXyvyilc40cXOKTkQ55EeYJwet1Sj1jtZWnRzIG32t0vgcjWRf
rmtCOMu4/fPeGU7Ba+LrCDm/+IDXnxPHqtG7l2+9kjlMRLfgpye/d/03QYS7BeLjEWfYEc9bS3VK
Mh43PW0Tbt8QRPx3nWd9JHeoFEbwY81XdXCFK2AnMHv+VVhM6d+U8RddyRomA0AZXie7HUP0sxz7
g1YCfouMpVXeD+GYx6DuEDVHAa85tkQ/u+3O9Ihs0tyLoCRSq0aTpZ8F8xUb/RCyR59xXgmDI793
FxN9b1gaPWeGqIkNLAdi8ZO088KSCwBTpPEuSsXTChd/bNxmWhHMfvu2tHtjo1idAT0Rn+6i/Ea9
OAqScSSFNbAcjnc5gJCB+f3Er9uz5rmOrE3leR0Z7vbLXtYl9z281KTjH2/mxFWhRQdWzJr9Fr2/
mgdWwmj+zwCdlf8nfKlhZiEiKMqBlWfjmsuaUnPzRiLXg0QN+bbJKOJO9YViyawtqr1d8I0PNVz4
iB/gosqsgD7XnVOjh3ZLkEYhNfk47rXk6iJzg7rIUoxDSz7KJsire5vqNFXcwj4G6q+oc26ORCmR
JbaKfZ7+NecnHTbl9BvrRRvL50WCQ85r7/JX1tUimZ2qsqPGGw4sh5eQnN7cLGJuQsAKqORR5AxP
tDGwbjZZSKx127QeQr2R68fViC12zF+lhA2TgmZg/7rknSKACguw3ftrayDIfDwwumIre2S02Df0
4rIJwFgJt1P8Qj96YnoVSgYd+5+0QtNO23Ee02IUSxamCRHUU3+vdfsgXnpuO4acow0CyARq2FZ4
5eyKb23b9WQllxOjYshIYQoyEUoYosQ+cYjh1NIBouqsSlSUySiBZCfEmpsujhl6QawwljR4ZLfF
ssGrJs29EeUmgmqFe+2/3/OHHb8Luyhw1EvxzbV2mE5ojDQmLBZZoZSOEheIkL9tOumifthNRrnQ
zWotsaa7qF/C8co1b3fDB2Pnyu78pEFmBK7EjsCCu9pgeWgWRqhWyQBQLZMaz3LyH0L7toiTTL7w
ZFrbdklCllb1ZJ1B/vst4a4D6VcKbqbHYmv8umZ4AENf0Oi5C8VpXBbgovMwbgorUdNPYibOlHTo
1Iv7fdcTlyvM2ssms3VARLTZB8lTBbjkfw+yIXtnF+ZJ9dSoYair0B4FaGKSglZ589nx3Cr3isls
dGSikfG5Qm+nHt2RjrjdhB/GGjssal99N1KA6p7VPn8hc8farhsAwxJi8s85kSZGnBmSf/6aFu+a
0jNeT9URKKG6aa235BuFdICpsHIUdfKMdTPNVALbuAZKhIQKcjrheFT5NJk7Z31BoeryJ5rPBb/B
pxWSv3qpvgkUkWRYmyY7DSjkm9N87Bhsku7aBJ0LRFOeN4wgI4NyeskRTsa5Y+JkfVkDJJaFcoNn
6906zvHwCRK46qWBwFkm4YY6DoucoESYMXojBCdThuPuYwsk5TKxokFBxtM1U92g/6OiUAGJV2ev
TiHIJUNmBN6wDjLxGDU0ndDYOP3uIQsCGbI/ZGyyw7WDsjtADcb5DXDBHJddfz4u/fn/ncRbQ1N4
1OxiTsM0fIdCDq9H4NG19RNppLlsMXs51HTHhDNnFKZLel+1BXhD6ozXlHiBtWW4Dp/Hjzx4by9R
46szgoq9HlRFdHitmsH33uHMb43pruJz8UoOys0Bd4dz3mL8LDkvcHT7zNw14lpT4KpgORXEFBEQ
hUiiHNuVOFQ+53zV36eSy3ZJtro6vPJFGzG8R41JipdtKqnukUwDO+6rsFkQd27yj7/vKiMTKcIq
znD+V7zRNSJTVJX/PlQvaZSEvZIsBIq/w0Hu/1z41zRaa88xnqHFV/q65cjkuMP5tvPxCfKfPSFS
A9L3dwiUdpL8FmtMAzvhu2FylX5lViC2bneMSXK8IbwSRx2qEe54vLB4Hf+O2YEvdit3K6BxkFkm
fGRgSTfHTgUYok/opuz8w6TXRWG451/xEJRcacnABI5i6m1yGXPMSXUDkBldB7NziJox9Q1zQWdb
K1dA1ryIfXiPHo8C82vkDKkM484noDK0FmNJCf30IPYsNRP3LUXiCPVovV9XBJoA0BKeHRfIIOCk
vqhiUDi5YhWhDvMU2c7zwkWK3BwBxsy9nN9CCNfQfbD7INTvuHUnYVRWgqrkN6L5+knuWumP/sPF
L6qY7ruGL2PZwCxkFtQFAoJ8ThWn6yBRfSfwdTxB9GOmKTUxT8sDeXo621qlBo60EdYJDxoFrKI5
gAoawo9bErKl3on+4bI8+93NsrjGgUegp6TGlkgvzXlii45lkxEiridvZNv1TtoX65CLRIUrYILj
ceAYwnMM1nwakEz9iVURmx5n/KP8MpSXdUg3B7GhuaA1AMCjBBVktJ7/IXIyoEX5AMuttCLEcJVo
aJeOLdkGgJJGkjnCuCiO69LqD2kJVCQkwmPw7my2tRit4Q4Vfp6NPnoqd01Sl9IMaR/2zjZDo+hD
ZYXegao2e5yGV6A8DY/bnEI+Ub/q2+W4qHXIBhjcfRFe+5Ipo8Fql2tZreLJszM6acT9AEm/nL+h
98ftnINiJZq3KLDCr4+AL919lbT2V7288Xr6C69kiwdqGbnqbRJ35OAs0hB0SLZn+iE+k5lZkUbC
HNiaU00XJe71q8bv+h5mzLw71HRkNzAt0ZsmL0Anb5h4nUN8RkmlyngONZjWh7r0rRs55bgmjQOU
X9ZrEyJj1IGES0phOJvKR7ZAegkpOelxcF1oe0ypk3+bUyklaSqexZevhu3ybTytd77MSfnXJkAg
dud2+Iv7c2ybgHrEJNrJj9c+A6cQp5JOuVvBigodXTw9O2imkRO9fD0zfa7SGdkbo6L5lbZH4ix8
KuNG+nwGzQOveePMgggHt8zc3fgdXtSdQyLkkpIV99CtqIYGURyGpbuxZDkLIHzshX3+LeDb3aR8
wwVSqkj8c+CNaHPA6xMPaoMyla5pejuKgHvdTMPRoYjUXZR22/rpsd7PpylEO1FJoqCs56y0Q9gQ
XAWmja/AvgkQHPcUfnuwSsWp4RUVrCVBc2nGMFWiXJB2DEw/mXaAUpmmZgk9/+JPHb0qh+Fw8MQR
JwQkpFTQOg9lHr1XXo6QmQFa3lQ8N1ooykOWvdFU28RmHqGzPSWsf8JySbUjVULpBMLJtUgFHy44
kVBhQytG4oZzYWHoXU3gR1vmljR3BfiFW6oSILUV/wpSLCyHsxHtJ+B9Uj5nh0FkNkRgRcj6rJUS
SZ3ATPKVVVxhfSd/+RiYJF8rJNegMaGKHnPslPaiAPNLZy2Cjrzw/uyIrrgFjpRfKnp8R3+fSVqp
S82Wy9L5JBhS9BHHgnYluwr0H0sZ/VeGAGjli99cdHrdLpLL9LhafgLHXdGaLJ9yq5GXrL7kV6mv
9UP/OFpzNvLwvfXHFMoQuWoiWdD2orQ+y2RRc1tzMeCxXWkHxYiCpYSaek8pLzaziXqQdezLW/RY
5naz6QqMpxi6cUy2u8itY2RBzTtTYVcYz9AEVIQSPuqoim16orz5DssYgE/vEMB/30ZAhJo7niLB
4ncsl5F+liAEMc3CsaGGJclZ6g3ioaZFJIEXyTBs+Qjdhd3sUOz5Ry9RP/LfuOmO1hKK98P03cnU
4E9UAZA6YIccw9qtwb/TyERc/cE//pfvreMr+C4AmVottrwzzkeQGimwWZ58C6OszO5Zqt4ARroV
PdgJaXkl+ATbyqBjTOTAI95KBUpzHYwL8OlIyk3yq4+TFYVo55yhiD1WSowu4faxKPgoN79Up/xj
d+psD8kwSdAc0kPA3EBWApAu29Q1OvtL0BHKVPXvR00g8wA9xhFKedC2SNHVuNsxR04KAuxUC7rz
fqctxTb8WcERzAp9JssjGFqUFaarAOTtxq3lqpprAf5yCxQts3oDS9LEWNWG4bzwSAZkZeY7L55w
ZogunlDMhdEUwBuAugnKu74+VTpE2MKiYOoiaCBkgF4d95qAj7iv8TmGijiW34pvyzJHSFLGRI1b
qNhLJHgVex4NHngACKx9vG4TQZg/wNRjJihcpMX5txHciFHzC+qJpDPMlgci1b9gD1uUmJZlAzcJ
piVmTTPiZqEftvWDIGX/Rbmie8oHLtLGzg6YiRWRj7/FWgbjJMPXhMKICfNnoyXHc/hvxPFn/p3J
JaAMGDyNEllewlnRJX/ffiBF2tw4E/CjciDLvWJwURKArJ3Jv6H4I+DPLVIjBgyI1ymTnPLABCXc
ytKV+nV0zvKwdWcU1LiSJ/YqVOip4N34Sk6nZhUj2BZ7H6B0+n93gBBK/YWfDvaNg0MQ5X2agBqw
hHtFyuGSL/R+4Z0jHIzeSVxYiblbx8nf0XdIpw3MsyFlmMgWL6s9yp2+mAmMn9LaE9qZhT/bTomD
wchpgU0Ggf8LH7YJmaxPBM26aY1iQjyX8GLWT7EZVWGFK6w4dgVGHSKRE78/gUoHSQ7UnomnR+eN
QPpkFhHBpgYEZLmwJbQ1ezoeCUD8XXTko2KQc7pYBGsmCDz0kSn0Dv7BbJmp1DMqXvLdcwA52PRh
uj3gd/bGAoptflKznc3Uf1xEgZsKxZ7JaVWkQ7Q7SLqa9KYV+l3S6Ve0JuOM6qoXxeFfMth+BmnR
bDM48AiwhgRiIes3xvNGM5YkOZuNFUnslosvR6N72SpRAPPOUnvHfTti2TPvzbuhFKAZ0N/+VnUp
dO21DJ7jc0gOMXYQnTNePgqd1kiORqIfeTrTPgb7wcQMYo9wCD1NOWNWhgPTC8h6q3qvxHKS88cu
OKYFmgH8yGX5qTmZR/0QvhWyATbjrs3oBK0QMDPpokrxrY+tMMVEZfx1po623xDG+GOvb/bwjF3i
zJZ/wCAj1es3z6BCB/OVzR3ExZqHCsb7fYW5Tke+HZJTGcp1TgEG7FQPOUPXyNXiY2cmDn8ZnMLG
DsH6i6o0zqbsB6v17U7Ey+Gpveorxb07tu0mdYWFqPUwNlgY5pLt/wg6vcj2Fka2P+kobbjeo6yV
vs2y9bQ4zKn6RktfWWMDfyWHKoZTYX7e+f1hwaTznKgvm0NjuRe3YF1bDTZQNiTci2vwDu0tnEpD
pz7TQdZoODPjphi2mAGgxK6S0TIX8O1t4Bze2kQE5IutW1KH5wuauKAwHHQQB+OdsJDunwX4cQv+
/aOqxlPidt8L+PSEtLLLUWAn7VvYdASMSQmKRQ4KUPJIaTBHXRTOfRmx/pj5QB1fWM3aeHR1HXwW
ZFcbT3if7XLLbeuxvMhjkDs5cgd6GBrRcyy/LP1jnlQ3g975JyJ7oBeVAjaSWPVji6o/nl5Z8vlP
FfHmsi7V6Bl6h/w6oQ7mTVXGd8+kC6K8YuNb+clVjTBVThVl74EIZp/h9vp3kFapSuvv/9AndO9H
RZcV0vtyNwLISKIMdXvRc99ovDi+4QDqANG2y5M0VPXdfh/IVicpJ9L41yR5Qt0P4p0uOZ/xbe+v
MaJl/9T8A2SfCREc6Gf1VLyrBEA1CbxJKoGUT3gUxXlYArn9mS9fo/QKQM0vDwEHJYMw5FGF3F89
ij4hE+rvqyhwCZzOarjvunj2KXmxl1OJFbOvglOJMADvn8qaV2YmaZFd2iMueLQuA1082QUVr/zF
cZdAcaGKr3/mSVqmII4Ax3YxRu4E4/18MB4RtrZq6RK2klv5TCMAYQmvMLAYc4kWznAIlkqY6MKT
D1F+A4WKOvN3SVujw6Lj6UHC0bQzMWqm951UN/oq8N50Hvtl4b8Y/PvkTIyyqa3z+SqjZbfczfI2
JlZ4yAhzjK+80KshCPj6uJqnv8Va9Vt1dWX3rgIjHto+VIDW9r4CrYibj5+0r2AVJoCQwINvnFMc
ioDsc1fV6FJqTi+xvVbH3WnM0wmB2WH42elCNtFAANGlciZF2rrYX1HSOifF6tC/cwd017wYziCq
13mC3bz8ooaqUvoYTtaBxh+afroOu0KtplNXJSvyjss527yKg/jfJV0iasDBln7R73ej8900Tn8o
qaM5nITawdcWsyqMOJbQCkE0XsosYegbYe3b18s2PvpmwMBKJcbiWxQ/gAn4gmrogp1pxsMhLvVh
7toeScvUTRTrp7zRpJSJKPPPGh19aWFduLMXHsieEA5Ry0zQn2/KrCZxpSRn7iWCyA45YIbKoT9j
iGYDHhgebnv2o3ogCMJAVdiKHmLIR9GDj4QMExeLMWpIVRwNXMgd+LccfSh/zfCcBGZGrrXkbZPE
jPmFY62cvu2qCTqZnJ2q32OCqiQy9hPxbBw73q87OB6BYEUwmU/ronN9Mr0fpXK8HcdhHUT4PsXa
cVHe1KVe9sDaZE2S8bpc2ETDTJImtTP9aVfw1G54Sc4EDlVlHjZCzlwN2p1LaauUT/I0sltaQPKY
cKwU/cfpGS+bJaW0dwYOvOGAWV8B+YgjUssmbUD9CmtEm7hFmWnbyIlQ13bsG83LU3f4PZ43kyjS
5gr7OkGyEyJUQYvLAveK6UfzXyDB94yEEWDuUTSC11qKnO+JFz+GnjGaGF7JzUz5naQsZZdhEz31
UrG4CXklIt+Nee3f5i/X/sO2Uhc/ERia86d2bs4LozbvW0jaK79y5/bIkVX47FwWvSjeMWkIaE7C
pWWp7v/RBWN6O8uSoPXLxODbZ5HKgsgnriPtWpAq1EtcFr8c58m9FZ0Fh0N0t1tPUR6LJDMd2psl
2lrnJ14VGJB7vqQG5wDgTmDfvw5szBFM6yGeP/O8GRQtjE5MPllPt5cc0RXycmQHd3X52Ff8XnXv
+MC9zvi7wb3+drnU8HrO43+OuDcKrOCI4FZcn38TKQfJP/cEIUsj02tOPv7knba8lK9Jl7e3fBsV
2OVpyl23JtYdFgJmk2/nCfoQPH+ni82Oj/DrsjSvSaQXU/vHiVflqPv3oElk9fkw04JGVjQ35Ytc
c3QfReMjNG93F00+A7fVG+8Il/Fp00FhWw/HAulTTXFbUdisnCvrs42ISfYNKTD69sFflirCq5c7
XGL5Zeju4oEmD7Vx5nEKD0fClInVbhFEMRZUrLpiN/dllHMRPXOmKpCics36lzxjddNPKr5IZ8Pk
jmWqCGU3rB43TGpx4FoeJ54+03BK0GMtOfCqcAzEyTvYC6ffsacD3yGqsRoSMi3NB2uD/PYUooXw
4KNdAIQhVrkzX4OVNN9tLgQI8lAMWkEuuVi559AW7lQbyU7TMoAKfcosO5xqtHe/a2zbMQ1Cj2eu
xPVheTujC3To3C+yswCmeof1W2GE744mCRMUmuI98J6psoDzDdrIlMcXgOyy7dViVwn5aYxZAeox
gGJnAW4cxlGUAXvu/zhIystt+DBIa9KOJ6SbXBIzt22dFHgb9KrT5T02h4H4QwGauX/XsV/lrdLk
nqveC77RFfuTuAGgEq9NUIn30yK0EkZFnWr7pfLLz0Vx4HnK+ohyHFJTCjqz1caZPdX5+mfpBonD
WAUDlZpR7GYQ7GTiZNDCExcsTsT7J2l3GtSR26bHUM3UdgGyqsWHZom2QGpPx+Ktbl9p6oIS5m1l
PdGURogI9vu3RRhYQSE5DGtoO2wp0y90T8+M7DWpzf011/37xjvp7chwe/XYf/R+lOWAzZmIqmZ2
wTMAY3oPbOCPM7xVrNdcFqagP2cc17NSTlOMIXANaV+jjnpWOs0GM6NgdqO6v/ZnKiBOLyWOe3EH
RhPnk8v0NyNvWVKOSw+xmdmCPyS7FftuBA17v2zQezWZoN7TgIgsbo9o1p394TO//HfronOvOMDm
v2XP4KHi8T321yfo3DyAHi6ZOhtLyJRBZK7X/2Xkt7p2gPuEMmMCtVTP+mUulmaDq2r+GoUF0gXt
m/QXMQXJWkmhCOsly1sWMbJ5Tgtu2whXI1/+nUDyY/c+8vCVF4H46b7aPollFtvuuvq5MJWfaj1R
ue9wyd5GxCyuzlTNP4KE7MAqK10e5jN5Ka+mBaPkSVSQEYwqWCIXxd/9kVQj76izruGnMW4w9XU7
SHGqDewb2zxOhNE5n/a8NwHI4tvY/KzarBCCjQuGseEZ5z2VMipnKe5xyHD2Oi7/GKJWjQmdHl8F
0uxxUKx+uWE5e5ryly/f71BiKlLh+9bYIHDtVfXnGqXU8OwONBr4OW1+LPCvYu079ilmtLHE+mjT
BqdMEmJ+FTtU8UhGGiLKRrXfOm+DV775FWZmeOmq28zWscSbnPK5hqwn27xqGpIhtMDxtOghcxTR
afhiHSoP8e6ayCfBtXHRLi55/XDHPSYm0IpcgVyPu8FjGaqP3KfOdVAHBHieJffxBkd0sV0MGYBY
yiRgDH6I6AX5b69XayZ1LIDvZmMDwOKPwpoNGWHT8eHURYKUehuUjWWjy1ooW2++IMia02+ujxS9
enwePCIUC44eRtImNHOhxuiyz79NSmh0GEA1hZckujtmyAulmt5aL4eYi4SXd8rAHWbI1/wKRWkN
Wvlf/nbOBzlle82bwpdIGDqkQiakokjXGIwf7sPquLUFJxBxXMPFgb8+DnHYUMjXXNbZYQjfkLEo
2nF+atWbLzh8TteEl+ysrlabBKAevx+BUYsxI2W0/skxuutM+n+1uTTUVoTC8L9ynPfZZXXbkWb1
cYbaSI8+q6TLYiRhtQTAKpwxaTrb/10rrYl7kRYU9T+KA9YobbhYPc/rHOZ3Kg5mwGEl0gJqCNB2
T1ZT14LbHmVdrBaz6+PT33hrIMV2/eP+HyFTjzkBIa2f/jchgx7qLSXbwkcgsvYJ5Hz0L1YiFXAU
8L7IgBtYr7BAPRKKv0ry4Yb/Tv177fk+KmKyXJ+v/v/+EPsoE6KiFXaefU5/dNbWLueiAjHoD+2N
uT57yTCVmiu/z99T3bTdOAlXxwIQSi5IzaB6MnKtPzq3bWiPbpL3b7MVI9kLmPxJ/flYgbCNC6nu
lA7Cl2sxYx8VEWG8RcvOwGup1yyeXFM8ZxpaNn+oOHLF9hApny4rj4u+DKpq+zzRJCkIBy73NtMk
s7IiM9G8Virp9IRTCcveET6pzHd40iX2m1zUb260E5HaGFUe/t3ueEi1+hXQdd725i1ZBrUXfHzG
t24/UTD1Gz5+6r5KOcWp3ZyYEKIHw0dpNNmKIqEJWTYbKwrJyedtSI08CVh+Q8c+5vCq2XRhjKrN
DLmtJksIOogp6iRrw3ecjtueQwGk/95mMMDpbWdkIXewrgz3iUAPzogHFGcZA5gOHuPM1H8IFsNa
B0ktYm8XLBS67yl/IG7Zj+tuBu/hpjU1GN85okYxZ5teDgHh/ANzLnDM/XvSOg1nDWD9x/KPFP+m
GDR/RM8MCrCie4tsBLA+Ly/JmjKrPmKvu0FAgdivlq2QUdpoRMtmqnTgtJJ73jWNoOlT7gRkMthX
lZddUeKqO9hJx9oHROz4JBcUPWDsucYYqy/F3qdbMFU32aYxgFI/dfeWrev/SweGPd2hSTCSWFS0
hBA71TP3ADvrOWyaNNjnIPFgTrPH3g2xYYvkpNDICURqz8ozap5AHJCU/o6Txpsd7XDyxmsX5WH7
6JGzqjuTa+8gHdprFue3UFlxlLOe59Ri3Ll7Q5OEub3DeF5CBFMjXtP/n3HdlglQ2QMUtJMJU9Cs
vQW8QjBPkpxUDn5n1D153ccz2zkXOlZtRpoylgMdpUq8fmT3+FzZk321Eg8TqlEdx+ZPF4gHL8zj
2Dhai5QNRgeLHygj6g1H7ZWL+imv1tkKHcHwgSGaC64s4FzAdThpByh8he/Xk5ZS//a/nIj2mZw1
bEFJTYSChobTCFO3FTp6W+uOTlQ/IXBRxn+YlbfhHX4eIYE6+wrFQjaUgletW0JXdP8j8QmDhg++
/DHss7vaZLqISV2nvLwGXBZ8b7cNneBGQyOqvxeeH2tODtqPWilOvroHBHVg2i/j+YxNJ9dGMy/z
FxxXb7DduQ9vZUWdGVkxgtoJZYqQVD3yxpIN8snBs3cQQwLwCzSY91h5P17j5n1SjPmR2cL5ILX5
CeUKRx4YtPXq8DnV8gym2R2gJaUrPHnTJ6FT+C2++FGyXqZ+mZoG23gvc1tdAsYcCAr8TW3unC6u
DMH09ikyk6+BA633Xz4aJFw/OOHQBMk4tWCDoxmuL47D4ofBcvBTqVDvzdwNOR/95vZEytB3UIek
55b0QYkzizZpDBkDQv3sU7DRQc/4Xxd3XY8wZ6TDADD376iRPJB06o2f8gwsU1XNa5LgIayGaNXc
7gcMeWliTUtNXam4nGNUbjnJtCyiUWKQmwNkWV0w9LsucjFabaQwsdjesGAcfftnguFBCFoyF7ae
OXok72YwSgxnJtm1YfOs5dmfCOhoc3x6NgmkfMUb/wqgmobqqIf80h761GSeHRy4D7680Qo67jGL
yvIQcQqexL0C0cMYPUIuAMkZRK/BQnqmKKmIT9xTkpn70oNoaZIK+EbVvgUt6gJID47aj1e7QCZW
UPC2OuD+QMJsLOudd6xOOVqiDaWXufKfe9eUfLxI9DEijsux08TP0PdLFOl4yZ34AHnLinlp8xmj
aLi8R13eFlwJp3aZGVP0kG0tOj82gu6xDF5PL7nfX0kBHApXeLiUPv3RVDEQwO4aZxJ2vKPhIb5s
Z7SblaP0GEcnK0rPzsBKmbKeCNhAxz6BI3G/Ps2xUq3K+F40YSGiHXcipN7w5yJdVjvQzWwdrxLS
Udpmw2YXLfsxu5gNyXiXIETAnzow71Jn4wEIHqRsam/xKqVdVSgOZgNbRzcDgZnsKPInTCIL4Ggi
yQjJ3GftUN39SoMXnp1z7F6TN28Iz/v+Pk/41QHAtOmLLLCWf2Py7mJPIXbDxOd0ncq4mifkXFLg
0M24yzlvt2y1ONBZyDgdvl6OFfMY7rB/Id3exMfUsGAkVQOhPCGuLDJwL/SrUeA4tEq6D6dhmIMM
llKXKpAkbLuN/S4d/uImJYArzJuWtZTbfEk8rFYzhX/McmIiQaSvuX4nZ+WUTE1g/qpCfj6S/ril
2DCKU0hEnYlviWFkng35iuNbDtQHAy/hPbIPWschM3uz3D8GygPBCxVsKt07/rcyRCEzhcqR4xB+
SxE41RtbKLimPHewaLTHDMBelpDsBW3h9IJvfu1yVYAVItrqD6BH5CsibssxfRoHXlDdjgwY2SkJ
HV2NbwLHmaB3CeB7HK1+h6wQfk8Epp6kwapxRsBVP8Dfiz5tKSoz3ugxFyHaIehnIMH6D+pvrZ8t
8cqZke09oXtCgxFQ7cD5QjQXcnVF8m17rqnI9tpoyiq503dcwhLoqqOg8tFO4BVcGyIYOUHCdAMY
WnZSXvK5UE7K7b3u8sFc3bPtQTatFqjJlaWnhrtfMQ4e8WKl5HUJK4bp2fVrPmkVW4qdBqiqNmeY
V/WXEVlO5Rm+9AehivTO0KK19AN+aTmd/JRYXMnqPZZ+YGFjqhNiOj0YFzhpWLI+BAlkg7S2CGdi
89vPN9I/WeC4C+hYUTnjCDPPd91Pq3h3h3kXNDlS/hj+2ZOpVQCP8CTuOC8yBj0IwGauC8LniLGu
rVMjSZH+P+mASFqnRTsYUBAkMk8ylCsLNXBFScHTVuC9VgyLIFuEWNC86cnq/hG8rb3MY0gNQkSf
lJp0j91UKWUqi+qHav4rjQI7+AF2jBY60c9xMZ7NHJbSs4P8qc/FwCRn+UnjC5/pSQF7OFUetCz4
aVM0SPl793/amw7Aocl1fYz4zvmjtGKEJ/HrvlE2oAxGkF6XmrsMdopqDsPe9XEQSUPekSLWKEHP
WHpcV3w+dRwxmgd1E4mHYkpP5pYBu7F3vWev9E3RNfTgaFV/bWCU1IszNHglIFoJP+JYAP0Yeo8F
k2Syd1eVvjKZSBU/L7MQMjF7R41udX+bXHBR2bjDSFLEW3PIZZIZplpoMalH/Xe1WQewR8/p7Dqs
2mC8WfgGXRiwz7jDEQSyzrUnE0FUWzaXixpjk6Gj4gEwapRBIA5WZwuv4DB6CtMicY20wiuFWov4
sslC2xTntT3yu+/ShQQNHPfzA3wDGqQhkdArOgJCbpESjleNil7lR/3ZZDGejpd2HqYApHnmI1i8
34tufLsTGrCJlUapxewJQddwbe9MuKasNbRZzFRtzTyiE+5jUR5s6FXCRNg0F3dZ52KZAWwecPHt
PlH2xaUfJsOLwvkfnwF4ipRlAux1hytlPRjxoXdqa1RJQmehe/hNJmVSq5w6R3xQ8TR2A1MU0ONg
Kwpt7OnEif0fj36wlhXDVm/LL1f44f6vlS8jfsMvsYNE6NRmMZF8jvB/LkSZPN4GOmZ9lLtz++Pm
z1kRaeEBTZSkSNGPCIhYSbiV7MHRvPVcQxIrMbq1d0IyYIW4o5tXwhI6G4kataG7ZZnX1XrivBMq
YsKxWDc0H95b43PzeOB2Fyb1Gw4hS7dDJucPll7DsZ7p2xRca9vyNT9Qvzc6XCYRcFWebDOspLRP
UCWR0P7pdbzW+/VqqioCpEWtHWZLVCjdoZzpY0MQh2NGvCVRuCj5sAWWV3mExH26U6EFN8D93Apc
7N793C6vdyPfWgETZvyhcfzIy0S/gEvAYkIoLYmwzLEwYpe23aYNcgE5k2vJk91AoGZ9LwvjHPpL
fMSkbuzxKaFoqFR7j8usnUrAKsM1do5G2cXWD4Rtr+GI596ajGhQPTi2UCG4sATiV+1QBX51dDwc
ZTcSO5eCKsGXlNtjL1mKPii7DCVJUjiexIxWTkCPLpTyaF2VNKzbXg/h351c4pPRSpUZwSeA57P8
YBay6SXcwPml7lgTEalD46fS0eQxJbb7pI/u9VA6nkejg/xWKi88S9iH4LfErJimSALxidPxyC+B
lGoIUJumemuX30zQxR2J+MNsdD8S/9xtqpXczbWBb5+SQUcZAVt9w6tHxZWEZH0lbFf5R2rmp4vF
eo7FbncnhBU3pnY5HLX4LQUaMOUq0x7a4wMcm32usVKIRadiZYnhhgsac00uyq3lR+KS+Z3N0LOq
2c+Vm7iSBzj3VeKsSUyuz+nv0YswHAEtdihNTOAtiplAEfDeGgOtdg9QEe9+LBp7Z9TUFWT84UCd
Qg0XRZTBpG5BSoBF1VI9CghCc7Ak4zU8GpPX5VUzPppzT54zPSr7/b954wsyiUELxjymOtx6GO96
qNL+hwfMvFGilMmzoilfwZGpmFqyMWbJPrjVOghrPxl5h0/LFCaxBXxYIueX0jXdWjtcZysZI9/U
AC6OYVcOLl/yDV+xcWCkqx6gwOU0Qtcznvm9OBiOZZIFBMzyNbqzbEMj2Ov8JeMIQwAo1pyDkSbr
dJBaQnwtQA9EV3GsUSIdrLO+DX70moEWGlqRnHNskduLwcxMmavzC+bz+xhV4f8b7dhj8j+zTB/w
gegh6eXUH01jehmmWEyNalgQygJy6dkh
`protect end_protected
